** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/OSC7.sch
.subckt OSC7 VDD VSS OUT_OSC7
*.PININFO VDD:B VSS:B OUT_OSC7:B
x8 VDD VSS net1 OUT_OSC7 inv_x4
x5 VDD VSS net2 net1 inv_x4
x6 VDD VSS net3 net2 inv_x4
x13 VDD VSS net4 net3 inv_x4
x14 VDD VSS net5 net4 inv_x4
x15 VDD VSS net6 net5 inv_x4
x16 VDD VSS OUT_OSC7 net6 inv_x4
.ends

* expanding   symbol:  inv_x4.sym # of pins=4
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/inv_x4.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/inv_x4.sch
.subckt inv_x4 VDD VSS INV_OUT INV_IN
*.PININFO INV_IN:I INV_OUT:O VDD:B VSS:B
XM3 INV_OUT INV_IN VDD VDD sky130_fd_pr__pfet_01v8 L=10 W=2 nf=1 m=1
XM5 INV_OUT INV_IN VSS VSS sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
.ends

.end
