magic
tech sky130A
timestamp 1770560933
<< error_s >>
rect 2000 1600 2028 1628
rect 4500 1600 4528 1628
rect 1972 1572 2000 1600
rect 4472 1572 4500 1600
rect 1972 -2100 2000 -2072
rect 4472 -2100 4500 -2072
rect 2000 -2128 2028 -2100
rect 4500 -2128 4528 -2100
<< metal1 >>
rect 6000 11100 6500 11200
rect 300 10800 800 10900
rect 2870 10800 5250 10810
rect 300 10500 5250 10800
rect 6000 10800 6100 11100
rect 6400 10800 6500 11100
rect 6000 10700 6500 10800
rect 7000 11100 7500 11200
rect 7000 10800 7100 11100
rect 7400 10800 7500 11100
rect 7000 10700 7500 10800
rect 8000 11100 8500 11200
rect 8000 10800 8100 11100
rect 8400 10800 8500 11100
rect 8000 10700 8500 10800
rect 9000 11100 9500 11200
rect 9000 10800 9100 11100
rect 9400 10800 9500 11100
rect 9000 10700 9500 10800
rect 10000 11100 10500 11200
rect 10000 10800 10100 11100
rect 10400 10800 10500 11100
rect 10000 10700 10500 10800
rect 11000 11100 11500 11200
rect 11000 10800 11100 11100
rect 11400 10800 11500 11100
rect 11000 10700 11500 10800
rect 12000 11100 12500 11200
rect 12000 10800 12100 11100
rect 12400 10800 12500 11100
rect 12000 10700 12500 10800
rect 13000 11100 13500 11200
rect 13000 10800 13100 11100
rect 13400 10800 13500 11100
rect 13000 10700 13500 10800
rect 300 10400 1000 10500
rect 2870 10400 12200 10500
rect 2870 10350 4500 10400
rect 2900 10300 3600 10350
rect 900 10090 1100 10100
rect 900 9810 910 10090
rect 1090 9810 1100 10090
rect 3100 10090 3300 10100
rect 900 9800 1100 9810
rect 1800 9850 2100 9900
rect 1800 9250 1850 9850
rect 2050 9250 2100 9850
rect 3100 9820 3110 10090
rect 3290 9820 3300 10090
rect 3100 9800 3300 9820
rect 4000 9950 4300 10000
rect 1800 9200 2100 9250
rect 3200 9200 3300 9300
rect 4000 9250 4050 9950
rect 4250 9250 4300 9950
rect 4000 9200 4300 9250
rect 800 9100 1000 9200
rect 600 8850 800 8900
rect 600 8750 650 8850
rect 750 8800 800 8850
rect 3150 8850 3350 8900
rect 750 8750 1000 8800
rect 600 8700 1000 8750
rect 3150 8750 3200 8850
rect 3300 8750 3350 8850
rect 5000 9800 12200 10400
rect 6700 9490 7900 9500
rect 6700 9410 6710 9490
rect 7030 9410 7900 9490
rect 6700 9400 7900 9410
rect 5400 9190 5700 9200
rect 5400 9110 5410 9190
rect 5690 9110 5700 9190
rect 5400 9100 5700 9110
rect 6760 9190 7750 9200
rect 6760 9110 6770 9190
rect 7090 9110 7750 9190
rect 6760 9100 7750 9110
rect 3150 8700 3350 8750
rect 5400 8500 5500 9100
rect 6750 8990 7600 9000
rect 6750 8910 6760 8990
rect 7080 8910 7600 8990
rect 6750 8900 7600 8910
rect 6760 8790 7450 8800
rect 6760 8710 6770 8790
rect 7090 8710 7450 8790
rect 6760 8700 7450 8710
rect 6760 8590 7300 8600
rect 6760 8510 6770 8590
rect 7090 8510 7300 8590
rect 7350 8550 7450 8700
rect 7500 8600 7600 8900
rect 7650 8750 7750 9100
rect 6760 8500 7300 8510
rect 3000 8490 3100 8500
rect 3090 8220 3100 8490
rect 5300 8300 5500 8500
rect 6750 8390 7100 8400
rect 6750 8310 6760 8390
rect 7080 8350 7100 8390
rect 7080 8310 7400 8350
rect 6750 8250 7400 8310
rect 3000 8200 3100 8220
rect 6760 8190 7550 8200
rect 6760 8110 6770 8190
rect 7090 8110 7550 8190
rect 6760 8100 7550 8110
rect 7600 8000 7700 8100
rect 6760 7990 7700 8000
rect 6760 7910 6770 7990
rect 7090 7910 7700 7990
rect 6760 7900 7700 7910
rect 2200 7400 2400 7500
rect 2700 7400 3500 7500
rect 0 7090 1150 7100
rect 0 6920 10 7090
rect 190 6920 1150 7090
rect 0 6900 1150 6920
rect 2200 6600 3500 7400
rect 10600 7000 13300 7800
rect 2200 6500 2400 6600
rect 2700 6500 3500 6600
rect 5900 6550 6150 6600
rect 5900 6350 5950 6550
rect 6100 6350 6150 6550
rect 11100 6400 11300 6500
rect 5900 6300 6150 6350
rect 12800 6200 13300 7000
rect 3000 6090 3200 6100
rect 3000 5810 3010 6090
rect 3190 5810 3200 6090
rect 11600 6000 13300 6200
rect 3000 5600 3200 5810
rect 5200 5780 5450 5800
rect 5200 5520 5270 5780
rect 5440 5520 5450 5780
rect 5200 5500 5450 5520
rect 11050 5550 11350 5600
rect 12100 5550 12700 5600
rect 600 5350 800 5400
rect 600 5250 650 5350
rect 750 5300 800 5350
rect 3200 5350 3400 5400
rect 750 5250 1000 5300
rect 600 5200 1000 5250
rect 3200 5250 3250 5350
rect 3350 5250 3400 5350
rect 11050 5350 11100 5550
rect 11300 5350 11350 5550
rect 12650 5350 12700 5550
rect 11050 5300 11350 5350
rect 12100 5300 12700 5350
rect 3200 5200 3400 5250
rect 900 4990 1100 5000
rect 900 4900 910 4990
rect 800 4800 910 4900
rect 900 4710 910 4800
rect 1090 4710 1100 4990
rect 3000 4800 3200 4900
rect 900 4700 1100 4710
rect 2800 4600 2900 4800
rect 4000 4750 4300 4800
rect 900 4190 1100 4200
rect 900 3910 910 4190
rect 1090 3910 1100 4190
rect 900 3900 1100 3910
rect 3100 4190 3300 4200
rect 3100 3910 3110 4190
rect 3290 3910 3300 4190
rect 3100 3900 3300 3910
rect 4000 3950 4050 4750
rect 4250 3950 4300 4750
rect 4000 3900 4300 3950
rect -300 3680 1300 3700
rect -300 3210 -290 3680
rect -110 3500 1300 3680
rect 1800 3500 2600 3600
rect 2900 3500 3500 3700
rect 4300 3500 4400 3700
rect -110 3400 1500 3500
rect 1800 3400 3900 3500
rect 4000 3400 4500 3500
rect -110 3210 1300 3400
rect 1800 3300 3500 3400
rect 4300 3300 4400 3400
rect -300 3200 1300 3210
rect 2600 3200 3700 3300
rect 1700 3100 2000 3200
rect 2600 2400 3500 3200
rect 5900 3850 6150 3900
rect 5900 3650 5950 3850
rect 6100 3650 6150 3850
rect 11200 3700 11300 3800
rect 5900 3600 6150 3650
rect 12800 3500 13300 6000
rect 5000 3400 5100 3500
rect 11600 3300 13300 3500
rect 11050 2850 11350 2900
rect 11050 2650 11100 2850
rect 11300 2650 11350 2850
rect 11050 2600 11350 2650
rect 12000 2850 12700 2900
rect 12000 2650 12050 2850
rect 12650 2650 12700 2850
rect 12000 2600 12700 2650
rect 2700 2090 2900 2100
rect 2700 1810 2710 2090
rect 2890 1810 2900 2090
rect 2700 1800 2900 1810
rect 5200 2090 5650 2100
rect 5200 1810 5430 2090
rect 5640 1810 5650 2090
rect 5200 1800 5650 1810
rect 900 1380 1100 1400
rect 900 1100 920 1380
rect 1090 1100 1100 1380
rect 900 1000 1100 1100
rect 600 750 1000 800
rect 600 650 650 750
rect 750 650 1000 750
rect 600 600 1000 650
rect 900 390 1100 400
rect 900 110 910 390
rect 1080 110 1100 390
rect 5900 1150 6150 1200
rect 3400 1000 3500 1100
rect 5900 950 5950 1150
rect 6100 950 6150 1150
rect 11000 1000 11400 1100
rect 5900 900 6150 950
rect 12800 800 13300 3300
rect 3100 750 3500 800
rect 3100 650 3150 750
rect 3250 650 3500 750
rect 3100 600 3500 650
rect 11600 600 13300 800
rect 3400 390 3600 400
rect 900 100 1100 110
rect 3400 110 3410 390
rect 3590 110 3600 390
rect 3400 100 3600 110
rect 4600 0 6600 600
rect 0 -110 1150 -100
rect 0 -390 10 -110
rect 190 -200 1150 -110
rect 1600 -200 3700 -100
rect 4400 -200 6600 0
rect 11050 150 11350 200
rect 11050 -50 11100 150
rect 11300 -50 11350 150
rect 11050 -100 11350 -50
rect 12000 150 12700 200
rect 12000 -50 12050 150
rect 12650 -50 12700 150
rect 12000 -100 12700 -50
rect 190 -300 1500 -200
rect 1600 -300 4100 -200
rect 4200 -300 6600 -200
rect 190 -390 1150 -300
rect 0 -400 1150 -390
rect 1700 -400 3700 -300
rect 4400 -500 6600 -300
rect 11000 -400 11400 -300
rect 900 -610 1100 -600
rect 900 -890 920 -610
rect 1090 -890 1100 -610
rect 3400 -610 3600 -600
rect 900 -900 1100 -890
rect 600 -1150 1100 -1100
rect 600 -1250 650 -1150
rect 750 -1250 1100 -1150
rect 600 -1300 1100 -1250
rect 900 -1600 1000 -1500
rect 3400 -890 3410 -610
rect 3590 -890 3600 -610
rect 3400 -900 3600 -890
rect 3100 -1150 3500 -1100
rect 3100 -1250 3150 -1150
rect 3250 -1250 3500 -1150
rect 4600 -1200 6600 -500
rect 3100 -1300 3500 -1250
rect 3400 -1600 3500 -1500
rect 5900 -1550 6150 -1500
rect 5900 -1750 5950 -1550
rect 6100 -1750 6150 -1550
rect 11000 -1700 11400 -1600
rect 5900 -1800 6150 -1750
rect 12800 -1900 13300 600
rect 11700 -2000 13300 -1900
rect 10900 -2100 13300 -2000
rect 10900 -2300 11700 -2100
rect 2700 -2350 3500 -2300
rect 2700 -2550 3200 -2350
rect 3450 -2550 3500 -2350
rect 2700 -2600 3500 -2550
rect 5200 -2310 5850 -2300
rect 5200 -2590 5710 -2310
rect 5840 -2590 5850 -2310
rect 5200 -2600 5850 -2590
rect 11050 -2550 11350 -2500
rect 11050 -2750 11100 -2550
rect 11300 -2750 11350 -2550
rect 11050 -2800 11350 -2750
rect 12000 -2550 12700 -2500
rect 12000 -2750 12050 -2550
rect 12650 -2750 12700 -2550
rect 12000 -2800 12700 -2750
rect -300 -3710 1200 -3700
rect -300 -3890 -290 -3710
rect -110 -3800 1200 -3710
rect 1300 -3800 4400 -3700
rect 5100 -3300 10900 -3000
rect 5100 -3500 5300 -3300
rect -110 -3890 4100 -3800
rect -300 -3900 4100 -3890
rect 5200 -4000 5600 -3900
rect 5200 -4200 5300 -4000
rect 5500 -4200 5600 -4000
rect 5200 -4300 5600 -4200
rect 7000 -4300 7200 -3300
rect 7300 -3850 7550 -3800
rect 7300 -4050 7350 -3850
rect 7500 -4050 7550 -3850
rect 7300 -4100 7550 -4050
rect 9000 -4300 9200 -3300
rect 9350 -3850 9600 -3800
rect 9350 -4050 9400 -3850
rect 9550 -4050 9600 -3850
rect 9350 -4100 9600 -4050
rect 11150 -3850 11400 -3800
rect 11150 -4050 11200 -3850
rect 11350 -4050 11400 -3850
rect 11150 -4100 11400 -4050
rect 12800 -4300 13300 -2100
rect 5800 -4500 13300 -4300
rect 9200 -4900 9500 -4850
rect 11050 -4900 11350 -4850
rect 5200 -4950 5500 -4900
rect 5200 -5150 5250 -4950
rect 5450 -5150 5500 -4950
rect 5200 -5200 5500 -5150
rect 6300 -4950 6900 -4900
rect 6300 -5150 6350 -4950
rect 6850 -5000 6900 -4950
rect 7200 -4950 7550 -4900
rect 6850 -5100 7000 -5000
rect 6850 -5150 6900 -5100
rect 6300 -5200 6900 -5150
rect 7200 -5150 7250 -4950
rect 7500 -5150 7550 -4950
rect 7200 -5200 7550 -5150
rect 8300 -4950 8900 -4900
rect 8300 -5150 8350 -4950
rect 8850 -5150 8900 -4950
rect 8300 -5200 8900 -5150
rect 9200 -5150 9250 -4900
rect 9450 -5150 9500 -4900
rect 9200 -5200 9500 -5150
rect 10300 -4950 10900 -4900
rect 10300 -5150 10350 -4950
rect 10850 -5150 10900 -4950
rect 10300 -5200 10900 -5150
rect 11050 -5150 11100 -4900
rect 11300 -5150 11350 -4900
rect 11050 -5200 11350 -5150
rect 12100 -4950 12700 -4900
rect 12100 -5150 12150 -4950
rect 12650 -5150 12700 -4950
rect 12100 -5200 12700 -5150
rect 12800 -5100 13300 -4500
rect 1800 -5500 1900 -5400
rect 2600 -5500 11900 -5400
rect 12800 -5500 13000 -5100
rect 1600 -5530 11900 -5500
rect 1600 -5880 1620 -5530
rect 2570 -5880 11900 -5530
rect 1600 -5900 11900 -5880
<< via1 >>
rect 6100 10800 6400 11100
rect 7100 10800 7400 11100
rect 8100 10800 8400 11100
rect 9100 10800 9400 11100
rect 10100 10800 10400 11100
rect 11100 10800 11400 11100
rect 12100 10800 12400 11100
rect 13100 10800 13400 11100
rect 910 9810 1090 10090
rect 1850 9250 2050 9850
rect 3110 9820 3290 10090
rect 4050 9250 4250 9950
rect 650 8750 750 8850
rect 3200 8750 3300 8850
rect 4500 8800 5000 10400
rect 6710 9410 7030 9490
rect 5410 9110 5690 9190
rect 6770 9110 7090 9190
rect 6760 8910 7080 8990
rect 6770 8710 7090 8790
rect 6770 8510 7090 8590
rect 2910 8220 3090 8490
rect 6760 8310 7080 8390
rect 6770 8110 7090 8190
rect 6770 7910 7090 7990
rect 2400 7400 2700 7700
rect 10 6920 190 7090
rect 2400 6300 2700 6600
rect 5950 6350 6100 6550
rect 3010 5810 3190 6090
rect 5270 5520 5440 5780
rect 650 5250 750 5350
rect 3250 5250 3350 5350
rect 11100 5350 11300 5550
rect 12050 5350 12650 5550
rect 910 4710 1090 4990
rect 910 3910 1090 4190
rect 3110 3910 3290 4190
rect 4050 3950 4250 4750
rect -290 3210 -110 3680
rect 4500 2400 5000 5200
rect 5950 3650 6100 3850
rect 11100 2650 11300 2850
rect 12050 2650 12650 2850
rect 2710 1810 2890 2090
rect 5430 1810 5640 2090
rect 920 1100 1090 1380
rect 650 650 750 750
rect 910 110 1080 390
rect 2100 200 2500 1300
rect 5950 950 6100 1150
rect 3150 650 3250 750
rect 3410 110 3590 390
rect 10 -390 190 -110
rect 11100 -50 11300 150
rect 12050 -50 12650 150
rect 920 -890 1090 -610
rect 650 -1250 750 -1150
rect 2100 -1800 2500 -700
rect 3410 -890 3590 -610
rect 3150 -1250 3250 -1150
rect 5950 -1750 6100 -1550
rect 3200 -2550 3450 -2350
rect 5710 -2590 5840 -2310
rect 11100 -2750 11300 -2550
rect 12050 -2750 12650 -2550
rect -290 -3890 -110 -3710
rect 4500 -3800 5000 -3000
rect 5300 -4200 5500 -4000
rect 7350 -4050 7500 -3850
rect 9400 -4050 9550 -3850
rect 11200 -4050 11350 -3850
rect 5250 -5150 5450 -4950
rect 6350 -5150 6850 -4950
rect 7250 -5150 7500 -4950
rect 8350 -5150 8850 -4950
rect 9250 -5150 9450 -4900
rect 10350 -5150 10850 -4950
rect 11100 -5150 11300 -4900
rect 12150 -5150 12650 -4950
rect 1620 -5880 2570 -5530
<< metal2 >>
rect 6000 11100 6500 11200
rect 6000 10800 6100 11100
rect 6400 10800 6500 11100
rect 400 10600 3300 10800
rect 6000 10700 6500 10800
rect 7000 11100 7500 11200
rect 7000 10800 7100 11100
rect 7400 10800 7500 11100
rect 7000 10700 7500 10800
rect 8000 11100 8500 11200
rect 8000 10800 8100 11100
rect 8400 10800 8500 11100
rect 8000 10700 8500 10800
rect 9000 11100 9500 11200
rect 9000 10800 9100 11100
rect 9400 10800 9500 11100
rect 9000 10700 9500 10800
rect 10000 11100 10500 11200
rect 10000 10800 10100 11100
rect 10400 10800 10500 11100
rect 10000 10700 10500 10800
rect 11000 11100 11500 11200
rect 11000 10800 11100 11100
rect 11400 10800 11500 11100
rect 11000 10700 11500 10800
rect 12000 11100 12500 11200
rect 12000 10800 12100 11100
rect 12400 10800 12500 11100
rect 12000 10700 12500 10800
rect 13000 11100 13500 11200
rect 13000 10800 13100 11100
rect 13400 10800 13500 11100
rect 13000 10700 13500 10800
rect 0 7090 200 7100
rect 0 6920 10 7090
rect 190 6920 200 7090
rect 0 6900 200 6920
rect -300 3680 -100 3700
rect -300 3210 -290 3680
rect -110 3210 -100 3680
rect -300 3200 -100 3210
rect 0 -110 200 -100
rect 0 -390 10 -110
rect 190 -390 200 -110
rect 0 -400 200 -390
rect 400 -3200 500 10600
rect 900 10090 1100 10600
rect 900 9810 910 10090
rect 1090 9810 1100 10090
rect 3100 10090 3300 10600
rect 600 8850 800 8900
rect 600 8750 650 8850
rect 750 8750 800 8850
rect 600 8700 800 8750
rect 600 5350 800 5400
rect 600 5250 650 5350
rect 750 5250 800 5350
rect 600 5200 800 5250
rect 900 4990 1100 9810
rect 1800 9850 2100 9900
rect 1800 9250 1850 9850
rect 2050 9250 2100 9850
rect 3100 9820 3110 10090
rect 3290 9820 3300 10090
rect 4400 10400 5100 10500
rect 3100 9800 3300 9820
rect 4000 9950 4300 10000
rect 1800 9200 2100 9250
rect 4000 9250 4050 9950
rect 4250 9250 4300 9950
rect 4000 9200 4300 9250
rect 3150 8850 3350 8900
rect 3150 8750 3200 8850
rect 3300 8750 3350 8850
rect 3150 8700 3350 8750
rect 4400 8800 4500 10400
rect 5000 8800 5100 10400
rect 5300 9650 5590 9680
rect 5300 9340 5320 9650
rect 5570 9500 5590 9650
rect 5570 9490 7100 9500
rect 5570 9410 6710 9490
rect 7030 9410 7100 9490
rect 5570 9400 7100 9410
rect 5570 9340 5590 9400
rect 5300 9310 5590 9340
rect 5400 9190 7100 9200
rect 5400 9110 5410 9190
rect 5690 9110 6770 9190
rect 7090 9110 7100 9190
rect 5400 9100 7100 9110
rect 2900 8490 3100 8500
rect 2900 8220 2910 8490
rect 3090 8220 3100 8490
rect 2900 8200 3100 8220
rect 2300 7700 2800 7800
rect 2300 7400 2400 7700
rect 2700 7400 2800 7700
rect 2300 7300 2800 7400
rect 2300 6600 2800 6700
rect 2300 6300 2400 6600
rect 2700 6300 2800 6600
rect 2300 6200 2800 6300
rect 3000 6090 3200 6100
rect 3000 5810 3010 6090
rect 3190 5810 3200 6090
rect 3000 5800 3200 5810
rect 3200 5350 3400 5400
rect 3200 5250 3250 5350
rect 3350 5250 3400 5350
rect 3200 5200 3400 5250
rect 4400 5200 5100 8800
rect 5300 8990 7100 9000
rect 5300 8910 6760 8990
rect 7080 8910 7100 8990
rect 5300 8900 7100 8910
rect 5300 6500 5350 8900
rect 5130 6480 5350 6500
rect 5130 6220 5140 6480
rect 5340 6220 5350 6480
rect 5130 6200 5350 6220
rect 5400 8790 7100 8800
rect 5400 8710 6770 8790
rect 7090 8710 7100 8790
rect 5400 8700 7100 8710
rect 5400 5800 5450 8700
rect 5250 5780 5450 5800
rect 5250 5520 5270 5780
rect 5440 5520 5450 5780
rect 5250 5500 5450 5520
rect 5500 8590 7100 8600
rect 5500 8510 6770 8590
rect 7090 8510 7100 8590
rect 5500 8500 7100 8510
rect 900 4710 910 4990
rect 1090 4710 1100 4990
rect 900 4190 1100 4710
rect 4000 4750 4300 4800
rect 900 3910 910 4190
rect 1090 3910 1100 4190
rect 900 3700 1100 3910
rect 3100 4190 3300 4200
rect 3100 3910 3110 4190
rect 3290 3910 3300 4190
rect 3100 3700 3300 3910
rect 4000 3950 4050 4750
rect 4250 3950 4300 4750
rect 4000 3900 4300 3950
rect 900 3400 3300 3700
rect 4400 2400 4500 5200
rect 5000 2400 5100 5200
rect 5500 3000 5550 8500
rect 5230 2990 5550 3000
rect 5230 2620 5250 2990
rect 5540 2620 5550 2990
rect 5230 2600 5550 2620
rect 5600 8390 7100 8400
rect 5600 8310 6760 8390
rect 7080 8310 7100 8390
rect 5600 8300 7100 8310
rect 12900 8300 13600 8700
rect 2700 2090 2900 2100
rect 2700 1810 2710 2090
rect 2890 1810 2900 2090
rect 2700 1800 2900 1810
rect 4400 1500 5100 2400
rect 5600 2100 5650 8300
rect 5420 2090 5650 2100
rect 5420 1810 5430 2090
rect 5640 1810 5650 2090
rect 5420 1800 5650 1810
rect 5700 8190 7100 8200
rect 5700 8110 6770 8190
rect 7090 8110 7100 8190
rect 5700 8100 7100 8110
rect 900 1380 1100 1400
rect 900 1100 920 1380
rect 1090 1100 1100 1380
rect 600 750 800 800
rect 600 650 650 750
rect 750 650 800 750
rect 600 600 800 650
rect 900 390 1100 1100
rect 2000 1300 2600 1400
rect 1700 700 1900 800
rect 900 110 910 390
rect 1080 110 1100 390
rect 900 -100 1100 110
rect 2000 200 2100 1300
rect 2500 200 2600 1300
rect 3500 1000 3700 1100
rect 3100 750 3300 800
rect 3100 650 3150 750
rect 3250 650 3300 750
rect 3100 600 3300 650
rect 2000 100 2600 200
rect 3400 390 3600 400
rect 3400 110 3410 390
rect 3590 110 3600 390
rect 4500 200 5100 1500
rect 3400 -100 3600 110
rect 900 -400 3600 -100
rect 900 -610 1100 -400
rect 900 -890 920 -610
rect 1090 -890 1100 -610
rect 900 -900 1100 -890
rect 2000 -700 2600 -600
rect 600 -1150 800 -1100
rect 600 -1250 650 -1150
rect 750 -1250 800 -1150
rect 600 -1300 800 -1250
rect 1700 -1300 1900 -1200
rect 2000 -1800 2100 -700
rect 2500 -1800 2600 -700
rect 2000 -1900 2600 -1800
rect -300 -3710 -100 -3700
rect -300 -3890 -290 -3710
rect -110 -3890 -100 -3710
rect -300 -3900 -100 -3890
rect 2900 -3900 3000 -400
rect 3400 -610 3600 -400
rect 3400 -890 3410 -610
rect 3590 -890 3600 -610
rect 3400 -900 3600 -890
rect 4400 -1000 5100 200
rect 3100 -1150 3300 -1100
rect 3100 -1250 3150 -1150
rect 3250 -1250 3300 -1150
rect 3100 -1300 3300 -1250
rect 3500 -1600 3700 -1500
rect 4500 -2000 5100 -1000
rect 5700 -1600 5750 8100
rect 5250 -1650 5750 -1600
rect 5250 -1850 5300 -1650
rect 5450 -1850 5750 -1650
rect 5250 -1900 5750 -1850
rect 5800 7990 7100 8000
rect 5800 7910 6770 7990
rect 7090 7910 7100 7990
rect 5800 7900 7100 7910
rect 3150 -2350 3500 -2300
rect 3150 -2550 3200 -2350
rect 3450 -2550 3500 -2350
rect 3150 -2600 3500 -2550
rect 4400 -3000 5100 -2000
rect 5800 -2300 5850 7900
rect 5900 6550 6150 6600
rect 5900 6350 5950 6550
rect 6100 6350 6150 6550
rect 5900 6300 6150 6350
rect 11050 5550 11350 5600
rect 11050 5350 11100 5550
rect 11300 5350 11350 5550
rect 11050 5300 11350 5350
rect 12000 5550 12700 5600
rect 12000 5350 12050 5550
rect 12650 5350 12700 5550
rect 12000 5300 12700 5350
rect 12800 5100 13600 8300
rect 11600 5000 13600 5100
rect 5900 3850 6150 3900
rect 5900 3650 5950 3850
rect 6100 3650 6150 3850
rect 5900 3600 6150 3650
rect 11050 2850 11350 2900
rect 11050 2650 11100 2850
rect 11300 2650 11350 2850
rect 11050 2600 11350 2650
rect 12000 2850 12700 2900
rect 12000 2650 12050 2850
rect 12650 2650 12700 2850
rect 12000 2600 12700 2650
rect 12800 2400 13600 5000
rect 11600 2300 13600 2400
rect 5900 1150 6150 1200
rect 5900 950 5950 1150
rect 6100 950 6150 1150
rect 5900 900 6150 950
rect 11050 150 11350 200
rect 11050 -50 11100 150
rect 11300 -50 11350 150
rect 11050 -100 11350 -50
rect 12000 150 12700 200
rect 12000 -50 12050 150
rect 12650 -50 12700 150
rect 12000 -100 12700 -50
rect 12800 -300 13600 2300
rect 11600 -400 13600 -300
rect 5900 -1550 6150 -1500
rect 5900 -1750 5950 -1550
rect 6100 -1750 6150 -1550
rect 5900 -1800 6150 -1750
rect 5700 -2310 5850 -2300
rect 5700 -2590 5710 -2310
rect 5840 -2590 5850 -2310
rect 5700 -2600 5850 -2590
rect 11050 -2550 11350 -2500
rect 11050 -2750 11100 -2550
rect 11300 -2750 11350 -2550
rect 11050 -2800 11350 -2750
rect 12000 -2550 12700 -2500
rect 12000 -2750 12050 -2550
rect 12650 -2750 12700 -2550
rect 12000 -2800 12700 -2750
rect 12800 -3000 13600 -400
rect 4400 -3800 4500 -3000
rect 5000 -3500 5100 -3000
rect 11600 -3100 13600 -3000
rect 4400 -3900 5000 -3800
rect 7300 -3850 7550 -3800
rect 5200 -4000 5600 -3900
rect 5200 -4200 5300 -4000
rect 5500 -4200 5600 -4000
rect 7300 -4050 7350 -3850
rect 7500 -4050 7550 -3850
rect 7300 -4100 7550 -4050
rect 9350 -3850 9600 -3800
rect 9350 -4050 9400 -3850
rect 9550 -4050 9600 -3850
rect 9350 -4100 9600 -4050
rect 11150 -3850 11400 -3800
rect 11150 -4050 11200 -3850
rect 11350 -4050 11400 -3850
rect 11150 -4100 11400 -4050
rect 12800 -3900 13600 -3100
rect 5200 -4300 5600 -4200
rect 9200 -4900 9500 -4850
rect 11050 -4900 11350 -4850
rect 5200 -4950 5500 -4900
rect 5200 -5150 5250 -4950
rect 5450 -5150 5500 -4950
rect 5200 -5200 5500 -5150
rect 6300 -4950 6900 -4900
rect 6300 -5150 6350 -4950
rect 6850 -5150 6900 -4950
rect 6300 -5200 6900 -5150
rect 7200 -4950 7550 -4900
rect 7200 -5150 7250 -4950
rect 7500 -5150 7550 -4950
rect 7200 -5200 7550 -5150
rect 8300 -4950 8900 -4900
rect 8300 -5150 8350 -4950
rect 8850 -5150 8900 -4950
rect 8300 -5200 8900 -5150
rect 9200 -5150 9250 -4900
rect 9450 -5150 9500 -4900
rect 9200 -5200 9500 -5150
rect 10300 -4950 10900 -4900
rect 10300 -5150 10350 -4950
rect 10850 -5150 10900 -4950
rect 10300 -5200 10900 -5150
rect 11050 -5150 11100 -4900
rect 11300 -5150 11350 -4900
rect 11050 -5200 11350 -5150
rect 12100 -4950 12700 -4900
rect 12100 -5150 12150 -4950
rect 12650 -5150 12700 -4950
rect 12100 -5200 12700 -5150
rect 12800 -5400 13000 -3900
rect 2200 -5500 13000 -5400
rect 1600 -5530 14100 -5500
rect 1600 -5880 1620 -5530
rect 2570 -5880 14100 -5530
rect 1600 -5900 14100 -5880
<< via2 >>
rect 6100 10800 6400 11100
rect 7100 10800 7400 11100
rect 8100 10800 8400 11100
rect 9100 10800 9400 11100
rect 10100 10800 10400 11100
rect 11100 10800 11400 11100
rect 12100 10800 12400 11100
rect 13100 10800 13400 11100
rect 10 6920 190 7090
rect -290 3210 -110 3680
rect 10 -390 190 -110
rect 650 8750 750 8850
rect 650 5250 750 5350
rect 1850 9250 2050 9850
rect 4050 9250 4250 9950
rect 3200 8750 3300 8850
rect 5320 9340 5570 9650
rect 2910 8220 3090 8490
rect 2400 7400 2700 7700
rect 2400 6300 2700 6600
rect 3010 5810 3190 6090
rect 3250 5250 3350 5350
rect 5140 6220 5340 6480
rect 4050 3950 4250 4750
rect 5250 2620 5540 2990
rect 2710 1810 2890 2090
rect 650 650 750 750
rect 2100 200 2500 1300
rect 3150 650 3250 750
rect 650 -1250 750 -1150
rect 2100 -1800 2500 -700
rect -290 -3890 -110 -3710
rect 3150 -1250 3250 -1150
rect 5300 -1850 5450 -1650
rect 3200 -2550 3450 -2350
rect 5950 6350 6100 6550
rect 11100 5350 11300 5550
rect 12050 5350 12650 5550
rect 5950 3650 6100 3850
rect 11100 2650 11300 2850
rect 12050 2650 12650 2850
rect 5950 950 6100 1150
rect 11100 -50 11300 150
rect 12050 -50 12650 150
rect 5950 -1750 6100 -1550
rect 11100 -2750 11300 -2550
rect 12050 -2750 12650 -2550
rect 5300 -4200 5500 -4000
rect 7350 -4050 7500 -3850
rect 9400 -4050 9550 -3850
rect 11200 -4050 11350 -3850
rect 5250 -5150 5450 -4950
rect 6350 -5150 6850 -4950
rect 7250 -5150 7500 -4950
rect 8350 -5150 8850 -4950
rect 9250 -5150 9450 -4900
rect 10350 -5150 10850 -4950
rect 11100 -5150 11300 -4900
rect 12150 -5150 12650 -4950
rect 1620 -5880 2570 -5530
<< metal3 >>
rect 6000 11100 6500 11200
rect 6000 10800 6100 11100
rect 6400 10800 6500 11100
rect 6000 10700 6500 10800
rect 7000 11100 7500 11200
rect 7000 10800 7100 11100
rect 7400 10800 7500 11100
rect 7000 10700 7500 10800
rect 8000 11100 8500 11200
rect 8000 10800 8100 11100
rect 8400 10800 8500 11100
rect 8000 10700 8500 10800
rect 9000 11100 9500 11200
rect 9000 10800 9100 11100
rect 9400 10800 9500 11100
rect 9000 10700 9500 10800
rect 10000 11100 10500 11200
rect 10000 10800 10100 11100
rect 10400 10800 10500 11100
rect 10000 10700 10500 10800
rect 11000 11100 11500 11200
rect 11000 10800 11100 11100
rect 11400 10800 11500 11100
rect 11000 10700 11500 10800
rect 12000 11100 12500 11200
rect 12000 10800 12100 11100
rect 12400 10800 12500 11100
rect 12000 10700 12500 10800
rect 13000 11100 13500 11200
rect 13000 10800 13100 11100
rect 13400 10800 13500 11100
rect 13000 10700 13500 10800
rect 600 10300 3400 10600
rect 600 8850 800 10300
rect 1800 9850 2100 9900
rect 1800 9250 1850 9850
rect 2050 9250 2100 9850
rect 1800 9200 2100 9250
rect 3200 9000 3400 10300
rect 4000 9950 4300 10000
rect 4000 9250 4050 9950
rect 4250 9250 4300 9950
rect 5300 9650 5590 9680
rect 5300 9340 5320 9650
rect 5570 9340 5590 9650
rect 5300 9310 5590 9340
rect 4000 9200 4300 9250
rect 600 8750 650 8850
rect 750 8750 800 8850
rect 600 7200 800 8750
rect 3150 8850 3400 9000
rect 3150 8750 3200 8850
rect 3300 8750 3400 8850
rect 3150 8700 3400 8750
rect 2900 8490 3100 8500
rect 2900 8210 2910 8490
rect 3090 8210 3100 8490
rect 2900 8200 3100 8210
rect 2300 7700 2800 7800
rect 2300 7400 2400 7700
rect 2700 7400 2800 7700
rect 2300 7300 2800 7400
rect 3200 7200 3400 8700
rect 0 7090 200 7100
rect 0 6920 10 7090
rect 190 6920 200 7090
rect 0 6900 200 6920
rect 600 6800 3400 7200
rect 600 5350 800 6800
rect 2300 6600 2800 6700
rect 2300 6300 2400 6600
rect 2700 6300 2800 6600
rect 2300 6200 2800 6300
rect 3000 6090 3200 6100
rect 3000 5810 3010 6090
rect 3190 5810 3200 6090
rect 3000 5800 3200 5810
rect 3300 5500 3400 6800
rect 5600 6550 6150 6600
rect 5130 6480 5350 6500
rect 5130 6220 5140 6480
rect 5340 6220 5350 6480
rect 5130 6200 5350 6220
rect 5600 6350 5950 6550
rect 6100 6350 6150 6550
rect 5600 6300 6150 6350
rect 600 5250 650 5350
rect 750 5250 800 5350
rect 600 3700 800 5250
rect 3100 5350 3400 5500
rect 3100 5250 3250 5350
rect 3350 5250 3400 5350
rect 3100 4500 3400 5250
rect 4000 4750 4300 4800
rect 3100 3700 3300 4500
rect 4000 3950 4050 4750
rect 4250 3950 4300 4750
rect 4000 3900 4300 3950
rect -300 3680 -100 3700
rect -300 3210 -290 3680
rect -110 3210 -100 3680
rect -300 3200 -100 3210
rect 600 3300 3300 3700
rect 600 750 800 3300
rect 2700 2090 2900 2100
rect 2700 1810 2710 2090
rect 2890 1810 2900 2090
rect 2700 1800 2900 1810
rect 600 650 650 750
rect 750 650 800 750
rect 600 -100 800 650
rect 2000 1300 2600 1400
rect 2000 200 2100 1300
rect 2500 200 2600 1300
rect 2000 100 2600 200
rect 3100 750 3300 3300
rect 5230 2990 5550 3000
rect 5230 2620 5250 2990
rect 5540 2620 5550 2990
rect 5230 2600 5550 2620
rect 3100 650 3150 750
rect 3250 650 3300 750
rect 3100 -100 3300 650
rect 0 -110 200 -100
rect 0 -390 10 -110
rect 190 -390 200 -110
rect 0 -400 200 -390
rect 600 -400 3300 -100
rect 600 -1150 800 -400
rect 600 -1250 650 -1150
rect 750 -1250 800 -1150
rect 600 -1400 800 -1250
rect 2000 -700 2600 -600
rect 2000 -1800 2100 -700
rect 2500 -1800 2600 -700
rect 3100 -1150 3300 -400
rect 3100 -1250 3150 -1150
rect 3250 -1250 3300 -1150
rect 3100 -1400 3300 -1250
rect 2000 -1900 2600 -1800
rect 5250 -1650 5500 -1600
rect 5250 -1850 5300 -1650
rect 5450 -1850 5500 -1650
rect 5250 -1900 5500 -1850
rect 3150 -2350 3500 -2300
rect 3150 -2550 3200 -2350
rect 3450 -2550 3500 -2350
rect 3150 -2600 3500 -2550
rect 5600 -3600 5650 6300
rect 11050 5550 11350 5600
rect 11050 5350 11100 5550
rect 11300 5350 11350 5550
rect 11050 5300 11350 5350
rect 12000 5550 12700 5600
rect 12000 5350 12050 5550
rect 12650 5350 12700 5550
rect 5200 -3700 5650 -3600
rect 5700 3850 6150 3900
rect 5700 3650 5950 3850
rect 6100 3650 6150 3850
rect 5700 3600 6150 3650
rect 5700 -3600 5750 3600
rect 11050 2850 11350 2900
rect 11050 2650 11100 2850
rect 11300 2650 11350 2850
rect 11050 2600 11350 2650
rect 12000 2850 12700 5350
rect 12000 2650 12050 2850
rect 12650 2650 12700 2850
rect 5800 1150 6150 1200
rect 5800 950 5950 1150
rect 6100 950 6150 1150
rect 5800 900 6150 950
rect 5800 -3450 5850 900
rect 11050 150 11350 200
rect 11050 -50 11100 150
rect 11300 -50 11350 150
rect 11050 -100 11350 -50
rect 12000 150 12700 2650
rect 12000 -50 12050 150
rect 12650 -50 12700 150
rect 5900 -1550 6150 -1500
rect 5900 -1750 5950 -1550
rect 6100 -1750 6150 -1550
rect 5900 -1800 6150 -1750
rect 5900 -3300 5950 -1800
rect 11050 -2550 11350 -2500
rect 11050 -2750 11100 -2550
rect 11300 -2750 11350 -2550
rect 11050 -2800 11350 -2750
rect 12000 -2550 12700 -50
rect 12000 -2750 12050 -2550
rect 12650 -2750 12700 -2550
rect 5900 -3400 11400 -3300
rect 5800 -3550 9600 -3450
rect 5700 -3700 7500 -3600
rect -300 -3710 -100 -3700
rect -300 -3890 -290 -3710
rect -110 -3890 -100 -3710
rect -300 -3900 -100 -3890
rect 5200 -4000 5600 -3700
rect 5200 -4200 5300 -4000
rect 5500 -4200 5600 -4000
rect 7300 -3800 7500 -3700
rect 7300 -3850 7550 -3800
rect 7300 -4050 7350 -3850
rect 7500 -4050 7550 -3850
rect 7300 -4100 7550 -4050
rect 9350 -3850 9600 -3550
rect 9350 -4050 9400 -3850
rect 9550 -4050 9600 -3850
rect 9350 -4100 9600 -4050
rect 11150 -3850 11400 -3400
rect 11150 -4050 11200 -3850
rect 11350 -4050 11400 -3850
rect 11150 -4100 11400 -4050
rect 5200 -4300 5600 -4200
rect 9200 -4900 9500 -4850
rect 11050 -4900 11350 -4850
rect 5200 -4950 5500 -4900
rect 5200 -5150 5250 -4950
rect 5450 -5150 5500 -4950
rect 5200 -5200 5500 -5150
rect 6300 -4950 6900 -4900
rect 6300 -5150 6350 -4950
rect 6850 -5150 6900 -4950
rect 6300 -5300 6900 -5150
rect 7200 -4950 7550 -4900
rect 7200 -5150 7250 -4950
rect 7500 -5150 7550 -4950
rect 7200 -5200 7550 -5150
rect 8300 -4950 8900 -4900
rect 8300 -5150 8350 -4950
rect 8850 -5150 8900 -4950
rect 8300 -5300 8900 -5150
rect 9200 -5150 9250 -4900
rect 9450 -5150 9500 -4900
rect 9200 -5200 9500 -5150
rect 10300 -4950 10900 -4900
rect 10300 -5150 10350 -4950
rect 10850 -5150 10900 -4950
rect 10300 -5300 10900 -5150
rect 11050 -5150 11100 -4900
rect 11300 -5150 11350 -4900
rect 11050 -5200 11350 -5150
rect 12000 -4950 12700 -2750
rect 12000 -5150 12150 -4950
rect 12650 -5150 12700 -4950
rect 12000 -5300 12700 -5150
rect 6300 -5500 12700 -5300
rect 1600 -5530 2600 -5500
rect 1600 -5880 1620 -5530
rect 2570 -5880 2600 -5530
rect 1600 -5900 2600 -5880
<< via3 >>
rect 6100 10800 6400 11100
rect 7100 10800 7400 11100
rect 8100 10800 8400 11100
rect 9100 10800 9400 11100
rect 10100 10800 10400 11100
rect 11100 10800 11400 11100
rect 12100 10800 12400 11100
rect 13100 10800 13400 11100
rect 1850 9250 2050 9850
rect 4050 9250 4250 9950
rect 5320 9340 5570 9650
rect 2910 8220 3090 8490
rect 2910 8210 3090 8220
rect 2400 7400 2700 7700
rect 10 6920 190 7090
rect 2400 6300 2700 6600
rect 3010 5810 3190 6090
rect 5140 6220 5340 6480
rect 4050 3950 4250 4750
rect -290 3210 -110 3680
rect 2710 1810 2890 2090
rect 2100 200 2500 1300
rect 5250 2620 5540 2990
rect 10 -390 190 -110
rect 2100 -1800 2500 -700
rect 5300 -1850 5450 -1650
rect 3200 -2550 3450 -2350
rect 11100 5350 11300 5550
rect 11100 2650 11300 2850
rect 11100 -50 11300 150
rect 11100 -2750 11300 -2550
rect -290 -3890 -110 -3710
rect 5250 -5150 5450 -4950
rect 7250 -5150 7500 -4950
rect 9250 -5150 9450 -4900
rect 11100 -5150 11300 -4900
rect 1620 -5880 2570 -5530
<< metal4 >>
rect 6000 11100 6500 11200
rect 300 10600 5900 10900
rect 0 7090 200 7200
rect 0 6920 10 7090
rect 190 6920 200 7090
rect 0 6800 200 6920
rect -300 3680 -100 3800
rect -300 3210 -290 3680
rect -110 3210 -100 3680
rect -300 3100 -100 3210
rect 0 -110 200 0
rect 0 -390 10 -110
rect 190 -390 200 -110
rect 0 -500 200 -390
rect 300 -3200 400 10600
rect 600 10300 4300 10500
rect 600 -3200 800 10300
rect 4000 9950 4300 10300
rect 900 9850 2100 9900
rect 900 9250 1850 9850
rect 2050 9250 2100 9850
rect 900 9200 2100 9250
rect 4000 9250 4050 9950
rect 4250 9250 4300 9950
rect 4000 9200 4300 9250
rect 5000 9650 5590 9690
rect 5000 9340 5320 9650
rect 5570 9340 5590 9650
rect 5000 9310 5590 9340
rect 5000 9200 5300 9310
rect 900 -3200 1100 9200
rect 4700 8900 5300 9200
rect 4700 8500 4900 8900
rect 2900 8490 4900 8500
rect 2900 8210 2910 8490
rect 3090 8210 4900 8490
rect 2900 8200 4900 8210
rect 2000 7700 2800 7800
rect 2000 7400 2400 7700
rect 2700 7400 2800 7700
rect 2000 6600 2800 7400
rect 2000 6300 2400 6600
rect 2700 6300 2800 6600
rect 2000 2900 2800 6300
rect 3000 6480 5350 6500
rect 3000 6220 5140 6480
rect 5340 6220 5350 6480
rect 3000 6200 5350 6220
rect 3000 6090 3200 6200
rect 3000 5810 3010 6090
rect 3190 5810 3200 6090
rect 3000 5800 3200 5810
rect 5700 4800 5900 10600
rect 4000 4750 5900 4800
rect 4000 3950 4050 4750
rect 4250 4300 5900 4750
rect 6000 10800 6100 11100
rect 6400 10800 6500 11100
rect 4250 3950 4300 4300
rect 4000 3900 4300 3950
rect 4600 2990 5550 3000
rect 2000 1300 2600 2900
rect 4600 2620 5250 2990
rect 5540 2620 5550 2990
rect 4600 2600 5550 2620
rect 4600 2100 4900 2600
rect 2700 2090 4900 2100
rect 2700 1810 2710 2090
rect 2890 1810 4900 2090
rect 2700 1800 4900 1810
rect 2000 200 2100 1300
rect 2500 200 2600 1300
rect 2000 100 2600 200
rect 2000 -700 2800 100
rect 2000 -1800 2100 -700
rect 2500 -1800 2800 -700
rect 2000 -1900 2800 -1800
rect 4600 -1650 5500 -1600
rect 4600 -1850 5300 -1650
rect 5450 -1850 5500 -1650
rect 4600 -1900 5500 -1850
rect 4600 -2300 4900 -1900
rect 3150 -2350 4900 -2300
rect 3150 -2550 3200 -2350
rect 3450 -2550 4900 -2350
rect 3150 -2600 4900 -2550
rect -300 -3710 -100 -3600
rect -300 -3890 -290 -3710
rect -110 -3890 -100 -3710
rect -300 -4000 -100 -3890
rect 6000 -4500 6500 10800
rect 5500 -4600 6500 -4500
rect 5148 -4950 6500 -4600
rect 5148 -5150 5250 -4950
rect 5450 -5150 6500 -4950
rect 5148 -5500 6500 -5150
rect 7000 11100 7500 11200
rect 7000 10800 7100 11100
rect 7400 10800 7500 11100
rect 7000 -4900 7500 10800
rect 8000 11100 8500 11200
rect 8000 10800 8100 11100
rect 8400 10800 8500 11100
rect 8000 -4500 8500 10800
rect 9000 11100 9500 11200
rect 9000 10800 9100 11100
rect 9400 10800 9500 11100
rect 9000 -3500 9500 10800
rect 10000 11100 10500 11200
rect 10000 10800 10100 11100
rect 10400 10800 10500 11100
rect 10000 -2000 10500 10800
rect 11000 11100 11500 11200
rect 11000 10800 11100 11100
rect 11400 10800 11500 11100
rect 11000 5550 11500 10800
rect 11000 5350 11100 5550
rect 11300 5350 11500 5550
rect 11000 5000 11500 5350
rect 12000 11100 12500 11200
rect 12000 10800 12100 11100
rect 12400 10800 12500 11100
rect 12000 3000 12500 10800
rect 11000 2850 12500 3000
rect 11000 2650 11100 2850
rect 11300 2650 12500 2850
rect 11000 2500 12500 2650
rect 13000 11100 13500 11200
rect 13000 10800 13100 11100
rect 13400 10800 13500 11100
rect 13000 500 13500 10800
rect 11000 150 13500 500
rect 11000 -50 11100 150
rect 11300 -50 13500 150
rect 11000 -500 13500 -50
rect 10000 -2550 11500 -2000
rect 10000 -2750 11100 -2550
rect 11300 -2750 11500 -2550
rect 10000 -3000 11500 -2750
rect 9000 -4000 11500 -3500
rect 8000 -4900 9500 -4500
rect 7000 -4950 7550 -4900
rect 7000 -5150 7250 -4950
rect 7500 -5150 7550 -4950
rect 7000 -5200 7550 -5150
rect 8000 -5150 9250 -4900
rect 9450 -5150 9500 -4900
rect 7000 -5500 7500 -5200
rect 8000 -5500 9500 -5150
rect 11000 -4900 11500 -4000
rect 11000 -5150 11100 -4900
rect 11300 -5150 11500 -4900
rect 11000 -5500 11500 -5150
rect 1600 -5530 2600 -5500
rect 1600 -5880 1620 -5530
rect 2570 -5880 2600 -5530
rect 1600 -5900 2600 -5880
use pdiscr  x0
timestamp 1770560933
transform 1 0 600 0 1 8500
box 400 -1500 2500 2000
use pdiscr  x1
timestamp 1770560933
transform 1 0 2800 0 1 8500
box 400 -1500 2500 2000
use pdiscr  x2
timestamp 1770560933
transform 1 0 600 0 -1 5500
box 400 -1500 2500 2000
use pdiscr  x3
timestamp 1770560933
transform 1 0 2800 0 -1 5500
box 400 -1500 2500 2000
use ndiscr  x4
timestamp 1770560933
transform 1 0 800 0 1 600
box 200 -800 2000 2800
use ndiscr  x5
timestamp 1770560933
transform 1 0 3300 0 1 600
box 200 -800 2000 2800
use ndiscr  x6
timestamp 1770560933
transform 1 0 800 0 -1 -1100
box 200 -800 2000 2800
use ndiscr  x7
timestamp 1770560933
transform 1 0 3300 0 -1 -1100
box 200 -800 2000 2800
use LOGIC  x8
timestamp 1770560933
transform 1 0 9100 0 1 8100
box -3100 -11100 4000 1900
use PASSGATE  x9
timestamp 1770560933
transform 1 0 11100 0 1 5800
box 200 -800 1619 911
use PASSGATE  x10
timestamp 1770560933
transform 1 0 11100 0 1 3100
box 200 -800 1619 911
use PASSGATE  x11
timestamp 1770560933
transform 1 0 11100 0 1 400
box 200 -800 1619 911
use PASSGATE  x12
timestamp 1770560933
transform 1 0 11100 0 1 -2300
box 200 -800 1619 911
use PASSGATE  x13
timestamp 1770560933
transform 1 0 5300 0 1 -4700
box 200 -800 1619 911
use PASSGATE  x14
timestamp 1770560933
transform 1 0 7300 0 1 -4700
box 200 -800 1619 911
use PASSGATE  x15
timestamp 1770560933
transform 1 0 9300 0 1 -4700
box 200 -800 1619 911
use PASSGATE  x16
timestamp 1770560933
transform 1 0 11100 0 1 -4700
box 200 -800 1619 911
<< labels >>
flabel metal1 900 8700 1000 8800 0 FreeSans 128 0 0 0 VCMUX_IN
port 20 nsew
flabel metal1 900 9100 1000 9200 0 FreeSans 128 0 0 0 vbg_0_2
port 19 nsew
flabel metal1 900 7000 1000 7100 0 FreeSans 128 0 0 0 VSS
port 13 nsew
flabel metal1 3200 9200 3300 9300 0 FreeSans 128 0 0 0 vbg_0_4
port 18 nsew
flabel metal1 900 4800 1000 4900 0 FreeSans 128 0 0 0 vbg_0_6
port 17 nsew
flabel metal1 3100 4800 3200 4900 0 FreeSans 128 0 0 0 vbg_0_8
port 16 nsew
flabel metal1 3400 1000 3500 1100 0 FreeSans 128 0 0 0 vbg_1_2
port 14 nsew
flabel metal1 900 1000 1000 1100 0 FreeSans 128 0 0 0 vbg_1_0
port 15 nsew
flabel metal1 900 -1600 1000 -1500 0 FreeSans 128 0 0 0 vbg_1_4
port 12 nsew
flabel metal1 3400 -1600 3500 -1500 0 FreeSans 128 0 0 0 vbg_1_6
port 10 nsew
flabel metal1 900 10400 1000 10500 0 FreeSans 128 0 0 0 VDD
port 11 nsew
flabel metal1 6400 11100 6500 11200 0 FreeSans 128 0 0 0 VCMUX_IN_1_0
port 4 nsew
flabel metal1 7400 11100 7500 11200 0 FreeSans 128 0 0 0 VCMUX_IN_1_2
port 3 nsew
flabel metal1 8400 11100 8500 11200 0 FreeSans 128 0 0 0 VCMUX_IN_1_4
port 2 nsew
flabel metal1 9400 11100 9500 11200 0 FreeSans 128 0 0 0 VCMUX_IN_1_6
port 0 nsew
flabel metal1 10400 11100 10500 11200 0 FreeSans 128 0 0 0 VCMUX_IN_0_8
port 5 nsew
flabel metal1 11400 11100 11500 11200 0 FreeSans 128 0 0 0 VCMUX_IN_0_2
port 8 nsew
flabel metal1 12400 11100 12500 11200 0 FreeSans 128 0 0 0 VCMUX_IN_0_4
port 7 nsew
flabel metal1 13400 11100 13500 11200 0 FreeSans 128 0 0 0 VCMUX_IN_0_6
port 6 nsew
flabel metal1 6900 -5100 7000 -5000 0 FreeSans 128 0 0 0 VCMUX_OUT
port 1 nsew
<< end >>
