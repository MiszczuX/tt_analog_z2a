magic
tech sky130A
timestamp 1769187801
<< metal1 >>
rect -2900 1700 -700 1800
rect -2900 -350 -2500 1700
rect -1400 1300 -800 1400
rect 3100 900 4000 1000
rect -1450 650 -1350 700
rect -1450 640 -1000 650
rect -1450 610 -1090 640
rect -1010 610 -1000 640
rect -1450 600 -1000 610
rect -1600 550 -1500 600
rect -1600 540 -900 550
rect -1600 510 -990 540
rect -910 510 -900 540
rect -1600 500 -900 510
rect -1750 450 -1650 500
rect -1750 440 -800 450
rect -1750 410 -890 440
rect -810 410 -800 440
rect -1750 400 -800 410
rect -1900 350 -1800 400
rect -1900 340 -700 350
rect -1900 310 -790 340
rect -710 310 -700 340
rect -1900 300 -700 310
rect -1800 240 -600 250
rect -1800 210 -690 240
rect -610 210 -600 240
rect -1800 200 -600 210
rect -1800 150 -1700 200
rect -1650 140 -500 150
rect -1650 110 -590 140
rect -510 110 -500 140
rect -1650 100 -500 110
rect 3900 100 4000 900
rect -1650 50 -1550 100
rect -1500 40 -430 50
rect -1500 10 -490 40
rect -440 10 -430 40
rect -1500 0 -430 10
rect 3500 0 4000 100
rect -1500 -50 -1400 0
rect -2900 -1075 -2850 -350
rect -2550 -1075 -2500 -350
rect -1500 -400 -1300 -300
rect -1200 -2660 -1150 -250
rect -1200 -2740 -1190 -2660
rect -1160 -2740 -1150 -2660
rect -1500 -3100 -1300 -2900
rect -1200 -3270 -1150 -2740
rect -1200 -3340 -1190 -3270
rect -1160 -3340 -1150 -3270
rect -1200 -8060 -1150 -3340
rect -1200 -8140 -1190 -8060
rect -1160 -8140 -1150 -8060
rect -1200 -8660 -1150 -8140
rect -1200 -8740 -1190 -8660
rect -1160 -8740 -1150 -8660
rect -2756 -10776 -2068 -10480
rect -2756 -11114 -2578 -10776
rect -2276 -10953 -2068 -10776
rect -1200 -10950 -1150 -8740
rect -1100 -2360 -1050 -250
rect -1100 -2440 -1090 -2360
rect -1060 -2440 -1050 -2360
rect -1100 -3560 -1050 -2440
rect -1100 -3630 -1090 -3560
rect -1060 -3630 -1050 -3560
rect -1100 -7760 -1050 -3630
rect -1100 -7840 -1090 -7760
rect -1060 -7840 -1050 -7760
rect -1100 -8960 -1050 -7840
rect -1100 -9040 -1090 -8960
rect -1060 -9040 -1050 -8960
rect -1100 -10950 -1050 -9040
rect -1000 -2060 -950 -250
rect -1000 -2140 -990 -2060
rect -960 -2140 -950 -2060
rect -1000 -3860 -950 -2140
rect -1000 -3940 -990 -3860
rect -960 -3940 -950 -3860
rect -1000 -7460 -950 -3940
rect -1000 -7540 -990 -7460
rect -960 -7540 -950 -7460
rect -1000 -9260 -950 -7540
rect -1000 -9340 -990 -9260
rect -960 -9340 -950 -9260
rect -1000 -10950 -950 -9340
rect -900 -1760 -850 -250
rect -900 -1840 -890 -1760
rect -860 -1840 -850 -1760
rect -900 -4160 -850 -1840
rect -900 -4240 -890 -4160
rect -860 -4240 -850 -4160
rect -900 -7160 -850 -4240
rect -900 -7240 -890 -7160
rect -860 -7240 -850 -7160
rect -900 -9560 -850 -7240
rect -900 -9640 -890 -9560
rect -860 -9640 -850 -9560
rect -900 -10950 -850 -9640
rect -800 -1460 -750 -250
rect -800 -1540 -790 -1460
rect -760 -1540 -750 -1460
rect -800 -4460 -750 -1540
rect -800 -4540 -790 -4460
rect -760 -4540 -750 -4460
rect -800 -6860 -750 -4540
rect -800 -6940 -790 -6860
rect -760 -6940 -750 -6860
rect -800 -10950 -750 -6940
rect -700 -4760 -650 -250
rect -700 -4840 -690 -4760
rect -660 -4840 -650 -4760
rect -700 -6560 -650 -4840
rect -700 -6640 -690 -6560
rect -660 -6640 -650 -6560
rect -700 -10950 -650 -6640
rect -600 -6260 -550 -250
rect -600 -6340 -590 -6260
rect -560 -6340 -550 -6260
rect -600 -10950 -550 -6340
rect -500 -10950 -450 -250
rect -400 -10950 -350 -100
rect -300 -2360 -250 -150
rect -300 -2440 -290 -2360
rect -260 -2440 -250 -2360
rect -300 -10950 -250 -2440
rect -200 -2060 -150 -150
rect -200 -2140 -190 -2060
rect -160 -2140 -150 -2060
rect -200 -3860 -150 -2140
rect -200 -3940 -190 -3860
rect -160 -3940 -150 -3860
rect -200 -10950 -150 -3940
rect -100 -1760 -50 -150
rect -100 -1840 -90 -1760
rect -60 -1840 -50 -1760
rect -100 -4160 -50 -1840
rect -100 -4240 -90 -4160
rect -60 -4240 -50 -4160
rect -100 -7160 -50 -4240
rect -100 -7240 -90 -7160
rect -60 -7240 -50 -7160
rect -100 -10950 -50 -7240
rect 0 -1460 50 -150
rect 0 -1540 10 -1460
rect 40 -1540 50 -1460
rect 0 -4460 50 -1540
rect 0 -4540 10 -4460
rect 40 -4540 50 -4460
rect 0 -6860 50 -4540
rect 0 -6940 10 -6860
rect 40 -6940 50 -6860
rect 0 -9860 50 -6940
rect 0 -9940 10 -9860
rect 40 -9940 50 -9860
rect 0 -10950 50 -9940
rect 100 -1160 150 -150
rect 100 -1240 110 -1160
rect 140 -1240 150 -1160
rect 100 -4760 150 -1240
rect 100 -4840 110 -4760
rect 140 -4840 150 -4760
rect 100 -6560 150 -4840
rect 100 -6640 110 -6560
rect 140 -6640 150 -6560
rect 100 -10160 150 -6640
rect 100 -10240 110 -10160
rect 140 -10240 150 -10160
rect 100 -10950 150 -10240
rect 200 -860 250 -150
rect 200 -940 210 -860
rect 240 -940 250 -860
rect 200 -3250 250 -940
rect 300 -560 350 -150
rect 500 -400 600 -300
rect 1600 -400 1800 -300
rect 300 -640 310 -560
rect 340 -640 350 -560
rect 200 -3350 240 -3250
rect 200 -5060 250 -3350
rect 200 -5140 210 -5060
rect 240 -5140 250 -5060
rect 200 -6260 250 -5140
rect 200 -6340 210 -6260
rect 240 -6340 250 -6260
rect 200 -10460 250 -6340
rect 200 -10540 210 -10460
rect 240 -10540 250 -10460
rect 200 -10950 250 -10540
rect 300 -5360 350 -640
rect 1900 -1700 2000 -1600
rect 400 -2450 500 -2400
rect 1800 -4000 1900 -2000
rect 2000 -4400 2100 -4300
rect 300 -5440 310 -5360
rect 340 -5440 350 -5360
rect 300 -5960 350 -5440
rect 300 -6040 310 -5960
rect 340 -6040 350 -5960
rect 300 -10760 350 -6040
rect 1900 -7100 2000 -7000
rect 500 -8500 600 -8400
rect 450 -8750 500 -8650
rect 450 -9050 550 -8950
rect 450 -9350 550 -9250
rect 1800 -7832 1900 -7400
rect 1800 -8832 3834 -7832
rect 1800 -9400 1900 -8832
rect 450 -9650 550 -9550
rect 1900 -9800 2000 -9700
rect 300 -10840 310 -10760
rect 340 -10840 350 -10760
rect 300 -10950 350 -10840
rect -2276 -11000 -1418 -10953
rect -2276 -11066 600 -11000
rect -2276 -11107 -1605 -11066
rect -1165 -11100 600 -11066
rect -2276 -11114 -2068 -11107
rect -2756 -11292 -2068 -11114
rect 2581 -11150 3393 -8832
rect -1569 -11205 -1278 -11165
rect 1968 -11205 5530 -11150
rect -1569 -11354 5530 -11205
rect -1569 -11357 2042 -11354
rect -1520 -11409 2042 -11357
<< via1 >>
rect -690 1310 -610 1390
rect -1090 610 -1010 640
rect -990 510 -910 540
rect -890 410 -810 440
rect -790 310 -710 340
rect -690 210 -610 240
rect -590 110 -510 140
rect 3500 100 3900 900
rect -490 10 -440 40
rect -2850 -1075 -2550 -350
rect -1190 -2740 -1160 -2660
rect -1190 -3340 -1160 -3270
rect -1190 -8140 -1160 -8060
rect -1190 -8740 -1160 -8660
rect -2578 -11114 -2276 -10776
rect -1090 -2440 -1060 -2360
rect -1090 -3630 -1060 -3560
rect -1090 -7840 -1060 -7760
rect -1090 -9040 -1060 -8960
rect -990 -2140 -960 -2060
rect -990 -3940 -960 -3860
rect -990 -7540 -960 -7460
rect -990 -9340 -960 -9260
rect -890 -1840 -860 -1760
rect -890 -4240 -860 -4160
rect -890 -7240 -860 -7160
rect -890 -9640 -860 -9560
rect -790 -1540 -760 -1460
rect -790 -4540 -760 -4460
rect -790 -6940 -760 -6860
rect -690 -4840 -660 -4760
rect -690 -6640 -660 -6560
rect -590 -6340 -560 -6260
rect -290 -2440 -260 -2360
rect -190 -2140 -160 -2060
rect -190 -3940 -160 -3860
rect -90 -1840 -60 -1760
rect -90 -4240 -60 -4160
rect -90 -7240 -60 -7160
rect 10 -1540 40 -1460
rect 10 -4540 40 -4460
rect 10 -6940 40 -6860
rect 10 -9940 40 -9860
rect 110 -1240 140 -1160
rect 110 -4840 140 -4760
rect 110 -6640 140 -6560
rect 110 -10240 140 -10160
rect 210 -940 240 -860
rect 310 -640 340 -560
rect 210 -5140 240 -5060
rect 210 -6340 240 -6260
rect 210 -10540 240 -10460
rect 1600 -3900 1800 -2100
rect 310 -5440 340 -5360
rect 310 -6040 340 -5960
rect 1600 -9300 1800 -7500
rect 310 -10840 340 -10760
<< metal2 >>
rect 3400 900 4000 1000
rect 3900 100 4000 900
rect -2587 -300 -1406 -255
rect -2900 -350 600 -300
rect -2900 -1075 -2850 -350
rect -2550 -400 600 -350
rect -2550 -442 -1406 -400
rect -2550 -765 -2500 -442
rect -1251 -560 700 -550
rect -1251 -640 310 -560
rect 340 -640 700 -560
rect -1251 -650 700 -640
rect -2550 -1075 -2482 -765
rect -1251 -860 700 -850
rect -1251 -940 210 -860
rect 240 -940 700 -860
rect -1251 -950 700 -940
rect -2733 -5443 -2482 -1075
rect -1251 -1160 700 -1150
rect -1251 -1240 110 -1160
rect 140 -1240 700 -1160
rect -1251 -1250 700 -1240
rect -1251 -1460 -750 -1450
rect -1251 -1540 -790 -1460
rect -760 -1540 -750 -1460
rect -1251 -1550 -750 -1540
rect 0 -1460 700 -1450
rect 0 -1540 10 -1460
rect 40 -1540 700 -1460
rect 0 -1550 700 -1540
rect -1251 -1760 -850 -1750
rect -1251 -1840 -890 -1760
rect -860 -1840 -850 -1760
rect -1251 -1850 -850 -1840
rect -100 -1760 700 -1750
rect -100 -1840 -90 -1760
rect -60 -1840 700 -1760
rect -100 -1850 700 -1840
rect 3500 -2000 4000 100
rect -1251 -2060 -950 -2050
rect -1251 -2140 -990 -2060
rect -960 -2140 -950 -2060
rect -1251 -2150 -950 -2140
rect -200 -2060 700 -2050
rect -200 -2140 -190 -2060
rect -160 -2140 700 -2060
rect -200 -2150 700 -2140
rect 1500 -2100 4000 -2000
rect -1251 -2360 -1050 -2350
rect -1251 -2440 -1090 -2360
rect -1060 -2440 -1050 -2360
rect -1251 -2450 -1050 -2440
rect -300 -2360 700 -2350
rect -300 -2440 -290 -2360
rect -260 -2440 700 -2360
rect -300 -2450 700 -2440
rect -1251 -2660 700 -2650
rect -1251 -2740 -1190 -2660
rect -1160 -2740 700 -2660
rect -1251 -2750 700 -2740
rect -1500 -3100 500 -2900
rect -1232 -3270 700 -3250
rect -1232 -3340 -1190 -3270
rect -1160 -3340 700 -3270
rect -1232 -3350 700 -3340
rect -1232 -3560 700 -3550
rect -1232 -3630 -1090 -3560
rect -1060 -3630 700 -3560
rect -1232 -3650 700 -3630
rect -1232 -3860 -950 -3850
rect -1232 -3940 -990 -3860
rect -960 -3940 -950 -3860
rect -1232 -3950 -950 -3940
rect -200 -3860 700 -3850
rect -200 -3940 -190 -3860
rect -160 -3940 700 -3860
rect -200 -3950 700 -3940
rect 1500 -3900 1600 -2100
rect 1800 -3000 4000 -2100
rect 1800 -3900 1900 -3000
rect 1500 -4000 1900 -3900
rect -1232 -4160 -850 -4150
rect -1232 -4240 -890 -4160
rect -860 -4240 -850 -4160
rect -1232 -4250 -850 -4240
rect -100 -4160 700 -4150
rect -100 -4240 -90 -4160
rect -60 -4240 700 -4160
rect -100 -4250 700 -4240
rect -1232 -4460 -750 -4450
rect -1232 -4540 -790 -4460
rect -760 -4540 -750 -4460
rect -1232 -4550 -750 -4540
rect 0 -4460 700 -4450
rect 0 -4540 10 -4460
rect 40 -4540 700 -4460
rect 0 -4550 700 -4540
rect -1232 -4760 -650 -4750
rect -1232 -4840 -690 -4760
rect -660 -4840 -650 -4760
rect -1232 -4850 -650 -4840
rect 100 -4760 700 -4750
rect 100 -4840 110 -4760
rect 140 -4840 700 -4760
rect 100 -4850 700 -4840
rect -1232 -5060 700 -5050
rect -1232 -5140 210 -5060
rect 240 -5140 700 -5060
rect -1232 -5150 700 -5140
rect -1232 -5360 700 -5350
rect -1232 -5440 310 -5360
rect 340 -5440 700 -5360
rect -2739 -5520 -2427 -5443
rect -1232 -5450 700 -5440
rect -2739 -5600 -1418 -5520
rect -2739 -5791 700 -5600
rect -2739 -10480 -2427 -5791
rect -1600 -5800 700 -5791
rect -1280 -5960 700 -5950
rect -1280 -6040 310 -5960
rect 340 -6040 700 -5960
rect -1280 -6050 700 -6040
rect -1280 -6260 -550 -6250
rect -1280 -6340 -590 -6260
rect -560 -6340 -550 -6260
rect -1280 -6350 -550 -6340
rect 200 -6260 700 -6250
rect 200 -6340 210 -6260
rect 240 -6340 700 -6260
rect 200 -6350 700 -6340
rect -1280 -6560 -650 -6550
rect -1280 -6640 -690 -6560
rect -660 -6640 -650 -6560
rect -1280 -6650 -650 -6640
rect 100 -6560 700 -6550
rect 100 -6640 110 -6560
rect 140 -6640 700 -6560
rect 100 -6650 700 -6640
rect -1280 -6860 -750 -6850
rect -1280 -6940 -790 -6860
rect -760 -6940 -750 -6860
rect -1280 -6950 -750 -6940
rect 0 -6860 700 -6850
rect 0 -6940 10 -6860
rect 40 -6940 700 -6860
rect 0 -6950 700 -6940
rect -1280 -7160 -850 -7150
rect -1280 -7240 -890 -7160
rect -860 -7240 -850 -7160
rect -1280 -7250 -850 -7240
rect -100 -7160 700 -7150
rect -100 -7240 -90 -7160
rect -60 -7240 700 -7160
rect -100 -7250 700 -7240
rect 1800 -7400 1900 -4000
rect -1280 -7460 700 -7450
rect -1280 -7540 -990 -7460
rect -960 -7540 700 -7460
rect -1280 -7550 700 -7540
rect 1500 -7500 1900 -7400
rect -1280 -7760 700 -7750
rect -1280 -7840 -1090 -7760
rect -1060 -7840 700 -7760
rect -1280 -7850 700 -7840
rect -1280 -8060 700 -8050
rect -1280 -8140 -1190 -8060
rect -1160 -8140 700 -8060
rect -1280 -8150 700 -8140
rect -1700 -8500 600 -8300
rect -1250 -8660 700 -8650
rect -1250 -8740 -1190 -8660
rect -1160 -8740 700 -8660
rect -1250 -8750 700 -8740
rect -1250 -8960 700 -8950
rect -1250 -9040 -1090 -8960
rect -1060 -9040 700 -8960
rect -1250 -9050 700 -9040
rect -1200 -9260 700 -9250
rect -1200 -9340 -990 -9260
rect -960 -9340 700 -9260
rect -1200 -9350 700 -9340
rect 1500 -9300 1600 -7500
rect 1800 -9300 1900 -7500
rect 1500 -9400 1900 -9300
rect -1250 -9560 700 -9550
rect -1250 -9640 -890 -9560
rect -860 -9640 700 -9560
rect -1250 -9650 700 -9640
rect -1200 -9860 700 -9850
rect -1200 -9940 10 -9860
rect 40 -9940 700 -9860
rect -1200 -9950 700 -9940
rect -1250 -10160 700 -10150
rect -1250 -10240 110 -10160
rect 140 -10240 700 -10160
rect -1250 -10250 700 -10240
rect -1300 -10460 700 -10450
rect -2756 -10776 -2068 -10480
rect -1300 -10540 210 -10460
rect 240 -10540 700 -10460
rect -1300 -10550 700 -10540
rect -2756 -11114 -2578 -10776
rect -2276 -11114 -2068 -10776
rect -1250 -10760 700 -10750
rect -1250 -10840 310 -10760
rect 340 -10840 700 -10760
rect -1250 -10850 700 -10840
rect -2756 -11292 -2068 -11114
use AND  x1
timestamp 1769186102
transform 1 0 450 0 1 -750
box 50 -2250 1550 450
use AND  x2
timestamp 1769186102
transform 1 0 450 0 -1 -5250
box 50 -2250 1550 450
use AND  x3
timestamp 1769186102
transform 1 0 450 0 1 -6150
box 50 -2250 1550 450
use AND  x4
timestamp 1769186102
transform 1 0 450 0 -1 -10650
box 50 -2250 1550 450
use LOGIC_INV  x9
timestamp 1769186102
transform 1 0 -1000 0 1 4600
box -200 -4850 4300 -2700
<< labels >>
flabel metal1 500 -8500 600 -8400 0 FreeSans 128 0 0 0 VSS
port 18 nsew
flabel metal1 500 -400 600 -300 0 FreeSans 128 0 0 0 VDD
port 17 nsew
flabel metal1 1900 -1700 2000 -1600 0 FreeSans 128 0 0 0 LOGICOUT_0_2
port 16 nsew
flabel metal1 1900 -7100 2000 -7000 0 FreeSans 128 0 0 0 LOGICOUT_0_6
port 14 nsew
flabel metal1 -1350 1300 -1250 1400 0 FreeSans 128 0 0 0 LOGICIN_0_2
port 12 nsew
flabel metal1 -1450 600 -1350 700 0 FreeSans 128 0 0 0 LOGICIN_0_4
port 11 nsew
flabel metal1 -1600 500 -1500 600 0 FreeSans 128 0 0 0 LOGICIN_0_6
port 10 nsew
flabel metal1 -1750 400 -1650 500 0 FreeSans 128 0 0 0 LOGICIN_0_8
port 8 nsew
flabel metal1 -1900 300 -1800 400 0 FreeSans 128 0 0 0 LOGICIN_1_0
port 7 nsew
flabel metal1 -1800 150 -1700 250 0 FreeSans 128 0 0 0 LOGICIN_1_2
port 6 nsew
flabel metal1 -1650 50 -1550 150 0 FreeSans 128 0 0 0 LOGICIN_1_4
port 5 nsew
flabel metal1 -1500 -50 -1400 50 0 FreeSans 128 0 0 0 LOGICIN_1_6
port 4 nsew
flabel metal1 2000 -4400 2100 -4300 0 FreeSans 128 0 0 0 LOGICOUT_0_4
port 15 nsew
rlabel metal1 -1569 -11357 -1363 -11205 1 VSS
port 18 n
flabel metal1 1900 -9800 2000 -9700 0 FreeSans 128 0 0 0 LOGICOUT_0_8
port 13 nsew
<< end >>
