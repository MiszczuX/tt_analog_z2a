magic
tech sky130A
magscale 1 2
timestamp 1770560933
<< viali >>
rect 1100 1740 2820 1800
rect 1040 820 1540 900
rect 1260 -100 1560 -40
rect 1260 -1400 1560 -1340
<< metal1 >>
rect 1080 1800 2840 1820
rect 1080 1680 1100 1800
rect 2820 1680 2840 1800
rect 1080 1660 2840 1680
rect 920 1400 980 1640
rect 1420 1520 1440 1580
rect 2700 1520 2720 1580
rect 1420 1500 2720 1520
rect 3060 1400 3120 1640
rect 400 1380 3200 1400
rect 400 1220 620 1380
rect 780 1220 3200 1380
rect 400 1200 3200 1220
rect 920 980 980 1200
rect 1400 1120 2980 1140
rect 1400 1060 1420 1120
rect 2700 1060 2980 1120
rect 3060 980 3120 1200
rect 1020 900 1600 960
rect 1020 820 1040 900
rect 1540 820 1600 900
rect 1020 200 1600 820
rect 400 0 1600 200
rect 1200 -40 1600 0
rect 1200 -100 1260 -40
rect 1560 -100 1600 -40
rect 1200 -120 1600 -100
rect 1800 -100 2600 0
rect 1800 -160 1900 -100
rect 1140 -200 1900 -160
rect 2500 -200 2600 -100
rect 1140 -220 2600 -200
rect 1180 -400 1380 -280
rect 800 -600 1380 -400
rect 400 -800 1380 -600
rect 800 -1000 1380 -800
rect 600 -1120 900 -1100
rect 600 -1280 620 -1120
rect 780 -1220 900 -1120
rect 1180 -1160 1380 -1000
rect 1440 -400 1620 -280
rect 1800 -300 2600 -220
rect 1440 -600 2000 -400
rect 1440 -800 3200 -600
rect 1440 -1000 2000 -800
rect 1440 -1160 1620 -1000
rect 780 -1280 1440 -1220
rect 600 -1300 900 -1280
rect 1200 -1340 1620 -1320
rect 1200 -1400 1260 -1340
rect 1560 -1400 1620 -1340
rect 400 -1420 1620 -1400
rect 400 -1580 1020 -1420
rect 1180 -1560 1620 -1420
rect 1180 -1580 1600 -1560
rect 400 -1600 1600 -1580
<< via1 >>
rect 1100 1740 2820 1760
rect 1100 1680 2820 1740
rect 1440 1520 2700 1580
rect 620 1220 780 1380
rect 1420 1060 2700 1120
rect 1900 -200 2500 -100
rect 620 -1280 780 -1120
rect 1020 -1580 1180 -1420
<< metal2 >>
rect 1000 1780 1200 1800
rect 1000 1760 2840 1780
rect 1000 1680 1100 1760
rect 2820 1680 2840 1760
rect 1000 1660 2840 1680
rect 600 1380 800 1400
rect 600 1220 620 1380
rect 780 1220 800 1380
rect 600 -1120 800 1220
rect 600 -1280 620 -1120
rect 780 -1280 800 -1120
rect 600 -1300 800 -1280
rect 1000 -1420 1200 1660
rect 1400 1520 1440 1580
rect 2700 1520 2720 1580
rect 1400 1120 2720 1520
rect 1400 1060 1420 1120
rect 2700 1060 2720 1120
rect 1800 -100 2600 1060
rect 1800 -200 1900 -100
rect 2500 -200 2600 -100
rect 1800 -300 2600 -200
rect 1000 -1580 1020 -1420
rect 1180 -1580 1200 -1420
rect 1000 -1600 1200 -1580
use sky130_fd_pr__nfet_01v8_64QSBY  sky130_fd_pr__nfet_01v8_64QSBY_0
timestamp 1770560933
transform 1 0 1411 0 1 -1121
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  sky130_fd_pr__pfet_01v8_MGS3BN_0
timestamp 1770560933
transform 1 0 1411 0 1 -316
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_A5ES5P  XM0pass
timestamp 1770560933
transform 0 1 2010 -1 0 1611
box -211 -1210 211 1210
use sky130_fd_pr__pfet_01v8_XGA8MR  XM1pass
timestamp 1770560933
transform 0 1 2019 -1 0 1011
box -211 -1219 211 1219
<< labels >>
flabel metal1 1000 -1600 1200 -1400 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 1000 0 1200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 800 -800 1000 -600 0 FreeSans 256 0 0 0 PASS_GATE_IN
port 1 nsew
flabel metal1 1800 -800 2000 -600 0 FreeSans 256 0 0 0 PASS_GATE_OUT
port 4 nsew
flabel metal1 400 1200 600 1400 0 FreeSans 256 0 0 0 PASS_GATE_EN
port 3 nsew
<< end >>
