magic
tech sky130A
magscale 1 2
timestamp 1765640399
<< checkpaint >>
rect 1035 -64 4849 42
rect 1035 -3098 7331 -64
rect 3517 -3204 7331 -3098
<< error_s >>
rect 2277 -1217 2312 -1200
rect 2278 -1218 2312 -1217
rect 2278 -1254 2348 -1218
rect 3536 -1254 3589 -1253
rect 2295 -1288 2366 -1254
rect 3518 -1288 3589 -1254
rect 4420 -1280 4460 -1255
rect 1586 -1320 1608 -1297
rect 1406 -1378 1430 -1362
rect 1402 -1488 1430 -1378
rect 1440 -1450 1480 -1328
rect 1492 -1378 1514 -1362
rect 1492 -1488 1518 -1378
rect 1240 -1613 1298 -1607
rect 1432 -1613 1490 -1607
rect 1624 -1613 1682 -1607
rect 1816 -1613 1874 -1607
rect 2008 -1613 2066 -1607
rect 1240 -1647 1252 -1613
rect 1432 -1647 1444 -1613
rect 1624 -1647 1636 -1613
rect 1816 -1647 1828 -1613
rect 2008 -1647 2020 -1613
rect 1240 -1653 1298 -1647
rect 1432 -1653 1490 -1647
rect 1624 -1653 1682 -1647
rect 1816 -1653 1874 -1647
rect 2008 -1653 2066 -1647
rect 2295 -1749 2365 -1288
rect 3519 -1289 3589 -1288
rect 2741 -1380 2760 -1322
rect 3536 -1323 3607 -1289
rect 4386 -1314 4494 -1289
rect 2769 -1356 2827 -1350
rect 2961 -1356 3019 -1350
rect 2769 -1390 2788 -1356
rect 2961 -1390 2973 -1356
rect 2577 -1396 2635 -1392
rect 2769 -1396 2827 -1390
rect 2961 -1396 3019 -1390
rect 3153 -1396 3211 -1392
rect 3345 -1396 3403 -1392
rect 2549 -1424 2663 -1420
rect 2741 -1424 2855 -1420
rect 2933 -1424 3047 -1420
rect 3125 -1424 3239 -1420
rect 3317 -1424 3431 -1420
rect 3226 -1440 3247 -1424
rect 2445 -1500 2671 -1440
rect 2445 -1616 2479 -1500
rect 2541 -1616 2575 -1500
rect 2637 -1616 2671 -1500
rect 3222 -1538 3247 -1440
rect 3260 -1500 3285 -1440
rect 3309 -1616 3343 -1440
rect 3405 -1616 3439 -1440
rect 2481 -1666 2539 -1660
rect 2673 -1666 2731 -1660
rect 2865 -1666 2923 -1660
rect 3057 -1666 3115 -1660
rect 3249 -1666 3307 -1660
rect 2481 -1700 2493 -1666
rect 2673 -1700 2685 -1666
rect 2865 -1700 2877 -1666
rect 3057 -1700 3069 -1666
rect 3249 -1700 3261 -1666
rect 2481 -1706 2539 -1700
rect 2673 -1706 2731 -1700
rect 2865 -1706 2923 -1700
rect 3057 -1706 3115 -1700
rect 3249 -1706 3307 -1700
rect 2295 -1785 2348 -1749
rect 3536 -1802 3606 -1323
rect 3790 -1380 3904 -1357
rect 3982 -1380 4096 -1357
rect 4174 -1380 4288 -1357
rect 3818 -1408 3876 -1385
rect 4010 -1408 4068 -1385
rect 4202 -1408 4260 -1385
rect 4394 -1391 4452 -1385
rect 4586 -1391 4644 -1385
rect 3818 -1425 3830 -1408
rect 4010 -1425 4022 -1408
rect 4202 -1425 4214 -1408
rect 4394 -1425 4406 -1391
rect 4586 -1425 4598 -1391
rect 3818 -1431 3876 -1425
rect 4010 -1431 4068 -1425
rect 4202 -1431 4260 -1425
rect 4394 -1431 4452 -1425
rect 4586 -1431 4644 -1425
rect 3722 -1719 3780 -1713
rect 3914 -1719 3972 -1713
rect 4106 -1719 4164 -1713
rect 4298 -1719 4356 -1713
rect 4490 -1719 4548 -1713
rect 3722 -1753 3734 -1719
rect 3914 -1753 3926 -1719
rect 4106 -1753 4118 -1719
rect 4298 -1753 4310 -1719
rect 4490 -1753 4502 -1719
rect 3722 -1759 3780 -1753
rect 3914 -1759 3972 -1753
rect 4106 -1759 4164 -1753
rect 4298 -1759 4356 -1753
rect 4490 -1759 4548 -1753
rect 3536 -1838 3589 -1802
<< viali >>
rect 1440 10 1480 200
rect 3480 180 3660 220
rect 1440 -1450 1480 -1270
rect 4420 -1280 4460 -1220
rect 2460 -1500 2660 -1440
rect 3260 -1500 3460 -1440
<< metal1 >>
rect 3450 240 3690 250
rect 1420 210 1490 220
rect 1420 200 1430 210
rect 1160 0 1430 200
rect 3450 160 3460 240
rect 3680 160 3690 240
rect 3450 150 3690 160
rect 1560 60 2760 120
rect 1420 -10 1490 0
rect 1530 10 1600 20
rect 1530 -50 1540 10
rect 1530 -60 1600 -50
rect 1720 10 1800 20
rect 1720 -50 1730 10
rect 1790 -50 1800 10
rect 1720 -60 1800 -50
rect 1910 10 1990 20
rect 1910 -50 1920 10
rect 1980 -50 1990 10
rect 1910 -60 1990 -50
rect 2100 10 2180 20
rect 2100 -50 2110 10
rect 2170 -50 2180 10
rect 2100 -60 2180 -50
rect 2290 10 2370 20
rect 2290 -50 2300 10
rect 2360 -50 2370 10
rect 2290 -60 2370 -50
rect 2490 10 2570 20
rect 2490 -50 2500 10
rect 2560 -50 2570 10
rect 2490 -60 2570 -50
rect 1620 -110 1700 -100
rect 1620 -170 1630 -110
rect 1690 -170 1700 -110
rect 1620 -180 1700 -170
rect 1810 -110 1890 -100
rect 1810 -170 1820 -110
rect 1880 -170 1890 -110
rect 1810 -180 1890 -170
rect 2004 -110 2080 -104
rect 2004 -170 2010 -110
rect 2070 -170 2080 -110
rect 2004 -176 2080 -170
rect 2200 -120 2280 -110
rect 2200 -180 2210 -120
rect 2270 -180 2280 -120
rect 1630 -190 1690 -180
rect 2200 -190 2280 -180
rect 2390 -120 2470 -110
rect 2390 -180 2400 -120
rect 2460 -180 2470 -120
rect 2390 -190 2470 -180
rect 2700 -220 2760 60
rect 1560 -280 2760 -220
rect 1580 -570 1700 -280
rect 1160 -770 1700 -570
rect 1580 -1000 1700 -770
rect 2700 -1000 2760 -280
rect 3150 60 4360 120
rect 3150 -220 3190 60
rect 3420 20 3500 30
rect 3420 -50 3430 20
rect 3490 -50 3500 20
rect 3420 -60 3500 -50
rect 3610 20 3690 30
rect 3610 -50 3620 20
rect 3680 -50 3690 20
rect 3610 -60 3690 -50
rect 3810 20 3890 30
rect 3810 -50 3820 20
rect 3880 -50 3890 20
rect 3810 -60 3890 -50
rect 4000 20 4080 30
rect 4000 -50 4010 20
rect 4070 -50 4080 20
rect 4000 -60 4080 -50
rect 4190 20 4270 30
rect 4190 -50 4200 20
rect 4260 -50 4270 20
rect 4190 -60 4270 -50
rect 3320 -100 3400 -90
rect 3320 -170 3330 -100
rect 3390 -170 3400 -100
rect 3320 -180 3400 -170
rect 3520 -100 3600 -90
rect 3520 -170 3530 -100
rect 3590 -170 3600 -100
rect 3520 -180 3600 -170
rect 3710 -100 3790 -90
rect 3710 -170 3720 -100
rect 3780 -170 3790 -100
rect 3710 -180 3790 -170
rect 3900 -100 3980 -90
rect 3900 -170 3910 -100
rect 3970 -170 3980 -100
rect 3900 -180 3980 -170
rect 4090 -100 4170 -90
rect 4090 -170 4100 -100
rect 4160 -170 4170 -100
rect 4090 -180 4170 -170
rect 4290 -100 4370 -90
rect 4290 -170 4300 -100
rect 4360 -170 4370 -100
rect 4290 -180 4370 -170
rect 3150 -280 4360 -220
rect 3150 -560 3190 -280
rect 2820 -570 3190 -560
rect 2820 -720 2830 -570
rect 2890 -720 3190 -570
rect 2820 -730 3190 -720
rect 1580 -1060 2760 -1000
rect 1620 -1100 1700 -1090
rect 1620 -1160 1630 -1100
rect 1690 -1160 1700 -1100
rect 1620 -1170 1700 -1160
rect 1810 -1100 1890 -1090
rect 1810 -1160 1820 -1100
rect 1880 -1160 1890 -1100
rect 1810 -1170 1890 -1160
rect 2010 -1100 2090 -1090
rect 2010 -1160 2020 -1100
rect 2080 -1160 2090 -1100
rect 2010 -1170 2090 -1160
rect 2200 -1100 2280 -1090
rect 2200 -1160 2210 -1100
rect 2270 -1160 2280 -1100
rect 2200 -1170 2280 -1160
rect 2390 -1100 2470 -1090
rect 2390 -1160 2400 -1100
rect 2460 -1160 2470 -1100
rect 2390 -1170 2470 -1160
rect 1430 -1220 1600 -1210
rect 1430 -1260 1530 -1220
rect 1160 -1270 1530 -1260
rect 1160 -1440 1400 -1270
rect 1510 -1280 1530 -1270
rect 1590 -1280 1600 -1220
rect 1510 -1290 1600 -1280
rect 1720 -1220 1800 -1210
rect 1720 -1280 1730 -1220
rect 1790 -1280 1800 -1220
rect 1720 -1290 1800 -1280
rect 1910 -1220 1990 -1210
rect 1910 -1280 1920 -1220
rect 1980 -1280 1990 -1220
rect 1910 -1290 1990 -1280
rect 2100 -1220 2180 -1210
rect 2100 -1280 2110 -1220
rect 2170 -1280 2180 -1220
rect 2100 -1290 2180 -1280
rect 2290 -1220 2370 -1210
rect 2290 -1280 2300 -1220
rect 2360 -1280 2370 -1220
rect 2290 -1290 2370 -1280
rect 2490 -1220 2570 -1210
rect 2490 -1280 2500 -1220
rect 2560 -1280 2570 -1220
rect 2490 -1290 2570 -1280
rect 1510 -1440 1530 -1290
rect 2700 -1320 2760 -1060
rect 1580 -1380 2760 -1320
rect 3150 -1000 3190 -730
rect 4480 -580 4830 -570
rect 4480 -760 4490 -580
rect 4550 -760 4830 -580
rect 4480 -770 4830 -760
rect 3150 -1060 4360 -1000
rect 3150 -1320 3190 -1060
rect 3420 -1100 3500 -1090
rect 3420 -1160 3430 -1100
rect 3490 -1160 3500 -1100
rect 3420 -1170 3500 -1160
rect 3620 -1100 3700 -1090
rect 3620 -1160 3630 -1100
rect 3690 -1160 3700 -1100
rect 3620 -1170 3700 -1160
rect 3810 -1100 3880 -1090
rect 3870 -1160 3880 -1100
rect 3810 -1170 3880 -1160
rect 4000 -1100 4080 -1090
rect 4000 -1160 4010 -1100
rect 4070 -1160 4080 -1100
rect 4000 -1170 4080 -1160
rect 4190 -1100 4270 -1090
rect 4190 -1160 4200 -1100
rect 4260 -1160 4270 -1100
rect 4190 -1170 4270 -1160
rect 4400 -1210 4480 -1200
rect 3320 -1220 3400 -1210
rect 3320 -1280 3330 -1220
rect 3390 -1280 3400 -1220
rect 3320 -1290 3400 -1280
rect 3520 -1220 3600 -1210
rect 3520 -1280 3530 -1220
rect 3590 -1280 3600 -1220
rect 3520 -1290 3600 -1280
rect 3710 -1220 3790 -1210
rect 3710 -1280 3720 -1220
rect 3780 -1280 3790 -1220
rect 3710 -1290 3790 -1280
rect 3900 -1220 3980 -1210
rect 3900 -1280 3910 -1220
rect 3970 -1280 3980 -1220
rect 3900 -1290 3980 -1280
rect 4090 -1220 4170 -1210
rect 4090 -1280 4100 -1220
rect 4160 -1280 4170 -1220
rect 4090 -1290 4170 -1280
rect 4290 -1220 4370 -1210
rect 4290 -1280 4300 -1220
rect 4360 -1280 4370 -1220
rect 4290 -1290 4370 -1280
rect 4400 -1290 4410 -1210
rect 4470 -1290 4480 -1210
rect 4400 -1300 4480 -1290
rect 3150 -1380 4360 -1320
rect 1160 -1450 1440 -1440
rect 1480 -1450 1530 -1440
rect 1160 -1460 1530 -1450
rect 2440 -1440 3560 -1420
rect 2440 -1500 2460 -1440
rect 2660 -1500 3260 -1440
rect 3460 -1500 3560 -1440
rect 2440 -1520 3560 -1500
<< via1 >>
rect 1430 200 1490 210
rect 1430 10 1440 200
rect 1440 10 1480 200
rect 1480 10 1490 200
rect 3460 220 3680 240
rect 3460 180 3480 220
rect 3480 180 3660 220
rect 3660 180 3680 220
rect 3460 160 3680 180
rect 1430 0 1490 10
rect 1540 -50 1600 10
rect 1730 -50 1790 10
rect 1920 -50 1980 10
rect 2110 -50 2170 10
rect 2300 -50 2360 10
rect 2500 -50 2560 10
rect 1630 -170 1690 -110
rect 1820 -170 1880 -110
rect 2010 -170 2070 -110
rect 2210 -180 2270 -120
rect 2400 -180 2460 -120
rect 3430 -50 3490 20
rect 3620 -50 3680 20
rect 3820 -50 3880 20
rect 4010 -50 4070 20
rect 4200 -50 4260 20
rect 3330 -170 3390 -100
rect 3530 -170 3590 -100
rect 3720 -170 3780 -100
rect 3910 -170 3970 -100
rect 4100 -170 4160 -100
rect 4300 -170 4360 -100
rect 2830 -720 2890 -570
rect 1630 -1160 1690 -1100
rect 1820 -1160 1880 -1100
rect 2020 -1160 2080 -1100
rect 2210 -1160 2270 -1100
rect 2400 -1160 2460 -1100
rect 1400 -1440 1440 -1270
rect 1440 -1440 1480 -1270
rect 1480 -1440 1510 -1270
rect 1530 -1280 1590 -1220
rect 1730 -1280 1790 -1220
rect 1920 -1280 1980 -1220
rect 2110 -1280 2170 -1220
rect 2300 -1280 2360 -1220
rect 2500 -1280 2560 -1220
rect 4490 -760 4550 -580
rect 3430 -1160 3490 -1100
rect 3630 -1160 3690 -1100
rect 3810 -1160 3870 -1100
rect 4010 -1160 4070 -1100
rect 4200 -1160 4260 -1100
rect 3330 -1280 3390 -1220
rect 3530 -1280 3590 -1220
rect 3720 -1280 3780 -1220
rect 3910 -1280 3970 -1220
rect 4100 -1280 4160 -1220
rect 4300 -1280 4360 -1220
rect 4410 -1220 4470 -1210
rect 4410 -1280 4420 -1220
rect 4420 -1280 4460 -1220
rect 4460 -1280 4470 -1220
rect 4410 -1290 4470 -1280
<< metal2 >>
rect 1370 210 1580 240
rect 1370 0 1430 210
rect 1490 20 1580 210
rect 3420 160 3460 240
rect 3680 160 3710 240
rect 3420 30 3710 160
rect 3420 20 4470 30
rect 1490 10 3430 20
rect 1490 0 1540 10
rect 1370 -50 1540 0
rect 1600 -50 1730 10
rect 1790 -50 1920 10
rect 1980 -50 2110 10
rect 2170 -50 2300 10
rect 2360 -50 2500 10
rect 2560 -50 3430 10
rect 3490 -50 3620 20
rect 3680 -50 3820 20
rect 3880 -50 4010 20
rect 4070 -50 4200 20
rect 4260 -50 4480 20
rect 1370 -60 4480 -50
rect 3320 -100 4550 -90
rect 1370 -110 2900 -100
rect 1370 -170 1630 -110
rect 1690 -170 1820 -110
rect 1880 -170 2010 -110
rect 2070 -120 2900 -110
rect 2070 -170 2210 -120
rect 1370 -180 2210 -170
rect 2270 -180 2400 -120
rect 2460 -180 2900 -120
rect 3320 -170 3330 -100
rect 3390 -170 3530 -100
rect 3590 -170 3720 -100
rect 3780 -170 3910 -100
rect 3970 -170 4100 -100
rect 4160 -170 4300 -100
rect 4360 -170 4550 -100
rect 3320 -180 4550 -170
rect 2200 -190 2280 -180
rect 2390 -190 2470 -180
rect 2822 -570 2898 -180
rect 2822 -720 2830 -570
rect 2890 -720 2898 -570
rect 1520 -1092 2570 -1090
rect 2822 -1092 2898 -720
rect 4480 -580 4550 -180
rect 4480 -760 4490 -580
rect 4480 -1090 4550 -760
rect 1520 -1100 2898 -1092
rect 1520 -1160 1630 -1100
rect 1690 -1160 1820 -1100
rect 1880 -1160 2020 -1100
rect 2080 -1160 2210 -1100
rect 2270 -1160 2400 -1100
rect 2460 -1160 2898 -1100
rect 1520 -1168 2898 -1160
rect 3320 -1100 4550 -1090
rect 3320 -1160 3430 -1100
rect 3490 -1160 3630 -1100
rect 3690 -1160 3810 -1100
rect 3870 -1160 4010 -1100
rect 4070 -1160 4200 -1100
rect 4260 -1160 4550 -1100
rect 1520 -1170 2570 -1168
rect 3320 -1170 4550 -1160
rect 1430 -1220 2570 -1210
rect 1430 -1260 1530 -1220
rect 1370 -1270 1530 -1260
rect 1370 -1440 1400 -1270
rect 1510 -1280 1530 -1270
rect 1590 -1280 1730 -1220
rect 1790 -1280 1920 -1220
rect 1980 -1280 2110 -1220
rect 2170 -1280 2300 -1220
rect 2360 -1280 2500 -1220
rect 2560 -1280 2570 -1220
rect 1510 -1290 2570 -1280
rect 3320 -1220 4410 -1210
rect 3320 -1280 3330 -1220
rect 3390 -1280 3530 -1220
rect 3590 -1280 3720 -1220
rect 3780 -1280 3910 -1220
rect 3970 -1280 4100 -1220
rect 4160 -1280 4300 -1220
rect 4360 -1280 4410 -1220
rect 3320 -1290 4410 -1280
rect 4470 -1290 4480 -1210
rect 1510 -1440 1610 -1290
rect 1370 -1460 1610 -1440
use sky130_fd_pr__pfet_01v8_8DVWZL  XM1
timestamp 1764261594
transform 1 0 1701 0 1 -1466
box -647 -319 647 319
use sky130_fd_pr__nfet_01v8_9DHFGX  XM2
timestamp 1764261594
transform 1 0 2942 0 1 -1528
box -647 -310 647 310
use sky130_fd_pr__pfet_01v8_8DVWZL  XM3
timestamp 1764261594
transform 1 0 4183 0 1 -1572
box -647 -319 647 319
use sky130_fd_pr__nfet_01v8_9DHFGX  XM4
timestamp 1764261594
transform 1 0 5424 0 1 -1634
box -647 -310 647 310
<< labels >>
flabel metal1 1160 0 1360 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 1160 -1460 1360 -1260 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 1160 -770 1360 -570 0 FreeSans 256 0 0 0 in_inv_amp
port 3 nsew
flabel metal1 4630 -770 4830 -570 0 FreeSans 256 0 0 0 out_amp_inv
port 2 nsew
<< end >>
