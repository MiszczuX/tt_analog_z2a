magic
tech sky130A
timestamp 1764263633
<< end >>
