magic
tech sky130A
timestamp 1769185602
<< metal1 >>
rect -2900 1700 -700 1800
rect -2900 -350 -2500 1700
rect -1400 1300 -800 1400
rect 3100 900 4000 1000
rect -1450 650 -1350 700
rect -1450 640 -1000 650
rect -1450 610 -1090 640
rect -1010 610 -1000 640
rect -1450 600 -1000 610
rect -1600 550 -1500 600
rect -1600 540 -900 550
rect -1600 510 -990 540
rect -910 510 -900 540
rect -1600 500 -900 510
rect -1750 450 -1650 500
rect -1750 440 -800 450
rect -1750 410 -890 440
rect -810 410 -800 440
rect -1750 400 -800 410
rect -1900 350 -1800 400
rect -1900 340 -700 350
rect -1900 310 -790 340
rect -710 310 -700 340
rect -1900 300 -700 310
rect -1800 240 -600 250
rect -1800 210 -690 240
rect -610 210 -600 240
rect -1800 200 -600 210
rect -1800 150 -1700 200
rect -1650 140 -500 150
rect -1650 110 -590 140
rect -510 110 -500 140
rect -1650 100 -500 110
rect 3900 100 4000 900
rect -1650 50 -1550 100
rect -1500 40 -430 50
rect -1500 10 -490 40
rect -440 10 -430 40
rect -1500 0 -430 10
rect 3500 0 4000 100
rect -1500 -50 -1400 0
rect -2900 -1097 -2850 -350
rect -2550 -1097 -2500 -350
rect -1500 -400 -1300 -300
rect -1500 -650 -1300 -550
rect -1500 -950 -1300 -850
rect -1500 -1250 -1300 -1150
rect -1500 -1550 -1300 -1450
rect -1500 -1850 -1300 -1750
rect -1500 -2150 -1300 -2050
rect -1500 -2450 -1300 -2350
rect -1500 -2750 -1300 -2650
rect -1200 -2660 -1150 -250
rect -1200 -2740 -1190 -2660
rect -1160 -2740 -1150 -2660
rect -1600 -2900 -1300 -2800
rect -1600 -3000 -1500 -2900
rect -1400 -3000 -1300 -2900
rect -1800 -3100 -1300 -3000
rect -1500 -3350 -1300 -3250
rect -1200 -3270 -1150 -2740
rect -1200 -3340 -1190 -3270
rect -1160 -3340 -1150 -3270
rect -1500 -3650 -1300 -3550
rect -1500 -3950 -1300 -3850
rect -1500 -4250 -1300 -4150
rect -1500 -4550 -1300 -4450
rect -1500 -4850 -1300 -4750
rect -1500 -5150 -1300 -5050
rect -1500 -5450 -1300 -5350
rect -1200 -5900 -1150 -3340
rect -1100 -2360 -1050 -250
rect -1100 -2440 -1090 -2360
rect -1060 -2440 -1050 -2360
rect -1100 -3560 -1050 -2440
rect -1100 -3630 -1090 -3560
rect -1060 -3630 -1050 -3560
rect -1100 -5900 -1050 -3630
rect -1000 -2060 -950 -250
rect -1000 -2140 -990 -2060
rect -960 -2140 -950 -2060
rect -1000 -3860 -950 -2140
rect -1000 -3940 -990 -3860
rect -960 -3940 -950 -3860
rect -1000 -5900 -950 -3940
rect -900 -1760 -850 -250
rect -900 -1840 -890 -1760
rect -860 -1840 -850 -1760
rect -900 -4160 -850 -1840
rect -900 -4240 -890 -4160
rect -860 -4240 -850 -4160
rect -900 -5900 -850 -4240
rect -800 -1460 -750 -250
rect -800 -1540 -790 -1460
rect -760 -1540 -750 -1460
rect -800 -4460 -750 -1540
rect -800 -4540 -790 -4460
rect -760 -4540 -750 -4460
rect -800 -5900 -750 -4540
rect -700 -4760 -650 -250
rect -700 -4840 -690 -4760
rect -660 -4840 -650 -4760
rect -700 -5900 -650 -4840
rect -600 -5900 -550 -250
rect -500 -5900 -450 -250
rect -400 -5900 -350 -100
rect -300 -2360 -250 -150
rect -300 -2440 -290 -2360
rect -260 -2440 -250 -2360
rect -300 -5900 -250 -2440
rect -200 -2060 -150 -150
rect -200 -2140 -190 -2060
rect -160 -2140 -150 -2060
rect -200 -3860 -150 -2140
rect -200 -3940 -190 -3860
rect -160 -3940 -150 -3860
rect -200 -5900 -150 -3940
rect -100 -1760 -50 -150
rect -100 -1840 -90 -1760
rect -60 -1840 -50 -1760
rect -100 -4160 -50 -1840
rect -100 -4240 -90 -4160
rect -60 -4240 -50 -4160
rect -100 -5900 -50 -4240
rect 0 -1460 50 -150
rect 0 -1540 10 -1460
rect 40 -1540 50 -1460
rect 0 -4460 50 -1540
rect 0 -4540 10 -4460
rect 40 -4540 50 -4460
rect 0 -5900 50 -4540
rect 100 -1160 150 -150
rect 100 -1240 110 -1160
rect 140 -1240 150 -1160
rect 100 -4760 150 -1240
rect 100 -4840 110 -4760
rect 140 -4840 150 -4760
rect 100 -5900 150 -4840
rect 200 -860 250 -150
rect 200 -940 210 -860
rect 240 -940 250 -860
rect 200 -3250 250 -940
rect 300 -560 350 -150
rect 500 -400 600 -300
rect 1600 -400 1800 -300
rect 300 -640 310 -560
rect 340 -640 350 -560
rect 200 -3350 240 -3250
rect 200 -5060 250 -3350
rect 200 -5140 210 -5060
rect 240 -5140 250 -5060
rect 200 -5900 250 -5140
rect 300 -5360 350 -640
rect 1900 -1700 2000 -1600
rect 400 -2450 500 -2400
rect 1800 -4000 1900 -2000
rect 2000 -4400 2100 -4300
rect 300 -5440 310 -5360
rect 340 -5440 350 -5360
rect 300 -5900 350 -5440
<< via1 >>
rect -690 1310 -610 1390
rect -1090 610 -1010 640
rect -990 510 -910 540
rect -890 410 -810 440
rect -790 310 -710 340
rect -690 210 -610 240
rect -590 110 -510 140
rect 3500 100 3900 900
rect -490 10 -440 40
rect -2850 -1097 -2550 -350
rect -1190 -2740 -1160 -2660
rect -1500 -3000 -1400 -2900
rect -1190 -3340 -1160 -3270
rect -1090 -2440 -1060 -2360
rect -1090 -3630 -1060 -3560
rect -990 -2140 -960 -2060
rect -990 -3940 -960 -3860
rect -890 -1840 -860 -1760
rect -890 -4240 -860 -4160
rect -790 -1540 -760 -1460
rect -790 -4540 -760 -4460
rect -690 -4840 -660 -4760
rect -290 -2440 -260 -2360
rect -190 -2140 -160 -2060
rect -190 -3940 -160 -3860
rect -90 -1840 -60 -1760
rect -90 -4240 -60 -4160
rect 10 -1540 40 -1460
rect 10 -4540 40 -4460
rect 110 -1240 140 -1160
rect 110 -4840 140 -4760
rect 210 -940 240 -860
rect 310 -640 340 -560
rect 210 -5140 240 -5060
rect 1600 -3900 1800 -2100
rect 310 -5440 340 -5360
<< metal2 >>
rect 3400 900 4000 1000
rect 3900 100 4000 900
rect -2900 -350 600 -300
rect -2900 -700 -2850 -350
rect -3100 -1097 -2850 -700
rect -2550 -400 600 -350
rect -2550 -700 -2500 -400
rect -1700 -560 700 -550
rect -1700 -640 310 -560
rect 340 -640 700 -560
rect -1700 -650 700 -640
rect -2550 -1097 -2400 -700
rect -1700 -860 700 -850
rect -1700 -940 210 -860
rect 240 -940 700 -860
rect -1700 -950 700 -940
rect -3100 -5600 -2400 -1097
rect -1700 -1160 700 -1150
rect -1700 -1240 110 -1160
rect 140 -1240 700 -1160
rect -1700 -1250 700 -1240
rect -1700 -1460 -750 -1450
rect -1700 -1540 -790 -1460
rect -760 -1540 -750 -1460
rect -1700 -1550 -750 -1540
rect 0 -1460 700 -1450
rect 0 -1540 10 -1460
rect 40 -1540 700 -1460
rect 0 -1550 700 -1540
rect -1700 -1760 -850 -1750
rect -1700 -1840 -890 -1760
rect -860 -1840 -850 -1760
rect -1700 -1850 -850 -1840
rect -100 -1760 700 -1750
rect -100 -1840 -90 -1760
rect -60 -1840 700 -1760
rect -100 -1850 700 -1840
rect 3500 -2000 4000 100
rect -1700 -2060 -950 -2050
rect -1700 -2140 -990 -2060
rect -960 -2140 -950 -2060
rect -1700 -2150 -950 -2140
rect -200 -2060 700 -2050
rect -200 -2140 -190 -2060
rect -160 -2140 700 -2060
rect -200 -2150 700 -2140
rect 1500 -2100 4000 -2000
rect -1700 -2360 -1050 -2350
rect -1700 -2440 -1090 -2360
rect -1060 -2440 -1050 -2360
rect -1700 -2450 -1050 -2440
rect -300 -2360 700 -2350
rect -300 -2440 -290 -2360
rect -260 -2440 700 -2360
rect -300 -2450 700 -2440
rect -1700 -2660 700 -2650
rect -1700 -2740 -1190 -2660
rect -1160 -2740 700 -2660
rect -1700 -2750 700 -2740
rect -1600 -2900 -1300 -2800
rect -1600 -3000 -1500 -2900
rect -1400 -3000 500 -2900
rect -1600 -3100 500 -3000
rect -1700 -3270 700 -3250
rect -1700 -3340 -1190 -3270
rect -1160 -3340 700 -3270
rect -1700 -3350 700 -3340
rect -1700 -3560 700 -3550
rect -1700 -3630 -1090 -3560
rect -1060 -3630 700 -3560
rect -1700 -3650 700 -3630
rect -1700 -3860 -950 -3850
rect -1700 -3940 -990 -3860
rect -960 -3940 -950 -3860
rect -1700 -3950 -950 -3940
rect -200 -3860 700 -3850
rect -200 -3940 -190 -3860
rect -160 -3940 700 -3860
rect -200 -3950 700 -3940
rect 1500 -3900 1600 -2100
rect 1800 -3000 4000 -2100
rect 1800 -3900 1900 -3000
rect 1500 -4000 1900 -3900
rect -1700 -4160 -850 -4150
rect -1700 -4240 -890 -4160
rect -860 -4240 -850 -4160
rect -1700 -4250 -850 -4240
rect -100 -4160 700 -4150
rect -100 -4240 -90 -4160
rect -60 -4240 700 -4160
rect -100 -4250 700 -4240
rect -1700 -4460 -750 -4450
rect -1700 -4540 -790 -4460
rect -760 -4540 -750 -4460
rect -1700 -4550 -750 -4540
rect 0 -4460 700 -4450
rect 0 -4540 10 -4460
rect 40 -4540 700 -4460
rect 0 -4550 700 -4540
rect -1700 -4760 -650 -4750
rect -1700 -4840 -690 -4760
rect -660 -4840 -650 -4760
rect -1700 -4850 -650 -4840
rect 100 -4760 700 -4750
rect 100 -4840 110 -4760
rect 140 -4840 700 -4760
rect 100 -4850 700 -4840
rect -1700 -5060 700 -5050
rect -1700 -5140 210 -5060
rect 240 -5140 700 -5060
rect -1700 -5150 700 -5140
rect -1700 -5360 700 -5350
rect -1700 -5440 310 -5360
rect 340 -5440 700 -5360
rect -1700 -5450 700 -5440
rect -3100 -5800 700 -5600
rect -3100 -5900 -1400 -5800
rect 1800 -6000 1900 -4000
use AND  x1
timestamp 1768672672
transform 1 0 450 0 1 -750
box 50 -2250 1550 450
use AND  x2
timestamp 1768672672
transform 1 0 450 0 -1 -5250
box 50 -2250 1550 450
use LOGIC_INV  x9
timestamp 1768674023
transform 1 0 -1000 0 1 4600
box -200 -4850 4300 -2700
<< labels >>
flabel metal1 500 -400 600 -300 0 FreeSans 128 0 0 0 VDD
port 17 nsew
flabel metal1 1900 -1700 2000 -1600 0 FreeSans 128 0 0 0 LOGICOUT_0_2
port 16 nsew
flabel metal1 -1350 1300 -1250 1400 0 FreeSans 128 0 0 0 LOGICIN_0_2
port 12 nsew
flabel metal1 -1450 600 -1350 700 0 FreeSans 128 0 0 0 LOGICIN_0_4
port 11 nsew
flabel metal1 -1600 500 -1500 600 0 FreeSans 128 0 0 0 LOGICIN_0_6
port 10 nsew
flabel metal1 -1750 400 -1650 500 0 FreeSans 128 0 0 0 LOGICIN_0_8
port 8 nsew
flabel metal1 -1900 300 -1800 400 0 FreeSans 128 0 0 0 LOGICIN_1_0
port 7 nsew
flabel metal1 -1800 150 -1700 250 0 FreeSans 128 0 0 0 LOGICIN_1_2
port 6 nsew
flabel metal1 -1650 50 -1550 150 0 FreeSans 128 0 0 0 LOGICIN_1_4
port 5 nsew
flabel metal1 -1500 -50 -1400 50 0 FreeSans 128 0 0 0 LOGICIN_1_6
port 4 nsew
flabel metal1 2000 -4400 2100 -4300 0 FreeSans 128 0 0 0 LOGICOUT_0_4
port 15 nsew
rlabel metal1 -1800 -3100 -1700 -3000 1 VSS
port 18 n
<< end >>
