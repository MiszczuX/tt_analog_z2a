magic
tech sky130A
magscale 1 2
timestamp 1768657996
<< nwell >>
rect -296 -1845 296 1845
<< pmos >>
rect -100 1426 100 1626
rect -100 990 100 1190
rect -100 554 100 754
rect -100 118 100 318
rect -100 -318 100 -118
rect -100 -754 100 -554
rect -100 -1190 100 -990
rect -100 -1626 100 -1426
<< pdiff >>
rect -158 1614 -100 1626
rect -158 1438 -146 1614
rect -112 1438 -100 1614
rect -158 1426 -100 1438
rect 100 1614 158 1626
rect 100 1438 112 1614
rect 146 1438 158 1614
rect 100 1426 158 1438
rect -158 1178 -100 1190
rect -158 1002 -146 1178
rect -112 1002 -100 1178
rect -158 990 -100 1002
rect 100 1178 158 1190
rect 100 1002 112 1178
rect 146 1002 158 1178
rect 100 990 158 1002
rect -158 742 -100 754
rect -158 566 -146 742
rect -112 566 -100 742
rect -158 554 -100 566
rect 100 742 158 754
rect 100 566 112 742
rect 146 566 158 742
rect 100 554 158 566
rect -158 306 -100 318
rect -158 130 -146 306
rect -112 130 -100 306
rect -158 118 -100 130
rect 100 306 158 318
rect 100 130 112 306
rect 146 130 158 306
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -306 -146 -130
rect -112 -306 -100 -130
rect -158 -318 -100 -306
rect 100 -130 158 -118
rect 100 -306 112 -130
rect 146 -306 158 -130
rect 100 -318 158 -306
rect -158 -566 -100 -554
rect -158 -742 -146 -566
rect -112 -742 -100 -566
rect -158 -754 -100 -742
rect 100 -566 158 -554
rect 100 -742 112 -566
rect 146 -742 158 -566
rect 100 -754 158 -742
rect -158 -1002 -100 -990
rect -158 -1178 -146 -1002
rect -112 -1178 -100 -1002
rect -158 -1190 -100 -1178
rect 100 -1002 158 -990
rect 100 -1178 112 -1002
rect 146 -1178 158 -1002
rect 100 -1190 158 -1178
rect -158 -1438 -100 -1426
rect -158 -1614 -146 -1438
rect -112 -1614 -100 -1438
rect -158 -1626 -100 -1614
rect 100 -1438 158 -1426
rect 100 -1614 112 -1438
rect 146 -1614 158 -1438
rect 100 -1626 158 -1614
<< pdiffc >>
rect -146 1438 -112 1614
rect 112 1438 146 1614
rect -146 1002 -112 1178
rect 112 1002 146 1178
rect -146 566 -112 742
rect 112 566 146 742
rect -146 130 -112 306
rect 112 130 146 306
rect -146 -306 -112 -130
rect 112 -306 146 -130
rect -146 -742 -112 -566
rect 112 -742 146 -566
rect -146 -1178 -112 -1002
rect 112 -1178 146 -1002
rect -146 -1614 -112 -1438
rect 112 -1614 146 -1438
<< nsubdiff >>
rect -260 1775 -164 1809
rect 164 1775 260 1809
rect -260 1713 -226 1775
rect 226 1713 260 1775
rect -260 -1775 -226 -1713
rect 226 -1775 260 -1713
rect -260 -1809 -164 -1775
rect 164 -1809 260 -1775
<< nsubdiffcont >>
rect -164 1775 164 1809
rect -260 -1713 -226 1713
rect 226 -1713 260 1713
rect -164 -1809 164 -1775
<< poly >>
rect -100 1707 100 1723
rect -100 1673 -84 1707
rect 84 1673 100 1707
rect -100 1626 100 1673
rect -100 1379 100 1426
rect -100 1345 -84 1379
rect 84 1345 100 1379
rect -100 1329 100 1345
rect -100 1271 100 1287
rect -100 1237 -84 1271
rect 84 1237 100 1271
rect -100 1190 100 1237
rect -100 943 100 990
rect -100 909 -84 943
rect 84 909 100 943
rect -100 893 100 909
rect -100 835 100 851
rect -100 801 -84 835
rect 84 801 100 835
rect -100 754 100 801
rect -100 507 100 554
rect -100 473 -84 507
rect 84 473 100 507
rect -100 457 100 473
rect -100 399 100 415
rect -100 365 -84 399
rect 84 365 100 399
rect -100 318 100 365
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -365 100 -318
rect -100 -399 -84 -365
rect 84 -399 100 -365
rect -100 -415 100 -399
rect -100 -473 100 -457
rect -100 -507 -84 -473
rect 84 -507 100 -473
rect -100 -554 100 -507
rect -100 -801 100 -754
rect -100 -835 -84 -801
rect 84 -835 100 -801
rect -100 -851 100 -835
rect -100 -909 100 -893
rect -100 -943 -84 -909
rect 84 -943 100 -909
rect -100 -990 100 -943
rect -100 -1237 100 -1190
rect -100 -1271 -84 -1237
rect 84 -1271 100 -1237
rect -100 -1287 100 -1271
rect -100 -1345 100 -1329
rect -100 -1379 -84 -1345
rect 84 -1379 100 -1345
rect -100 -1426 100 -1379
rect -100 -1673 100 -1626
rect -100 -1707 -84 -1673
rect 84 -1707 100 -1673
rect -100 -1723 100 -1707
<< polycont >>
rect -84 1673 84 1707
rect -84 1345 84 1379
rect -84 1237 84 1271
rect -84 909 84 943
rect -84 801 84 835
rect -84 473 84 507
rect -84 365 84 399
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -399 84 -365
rect -84 -507 84 -473
rect -84 -835 84 -801
rect -84 -943 84 -909
rect -84 -1271 84 -1237
rect -84 -1379 84 -1345
rect -84 -1707 84 -1673
<< locali >>
rect -260 1775 -164 1809
rect 164 1775 260 1809
rect -260 1713 -226 1775
rect 226 1713 260 1775
rect -100 1673 -84 1707
rect 84 1673 100 1707
rect -146 1614 -112 1630
rect -146 1422 -112 1438
rect 112 1614 146 1630
rect 112 1422 146 1438
rect -100 1345 -84 1379
rect 84 1345 100 1379
rect -100 1237 -84 1271
rect 84 1237 100 1271
rect -146 1178 -112 1194
rect -146 986 -112 1002
rect 112 1178 146 1194
rect 112 986 146 1002
rect -100 909 -84 943
rect 84 909 100 943
rect -100 801 -84 835
rect 84 801 100 835
rect -146 742 -112 758
rect -146 550 -112 566
rect 112 742 146 758
rect 112 550 146 566
rect -100 473 -84 507
rect 84 473 100 507
rect -100 365 -84 399
rect 84 365 100 399
rect -146 306 -112 322
rect -146 114 -112 130
rect 112 306 146 322
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -322 -112 -306
rect 112 -130 146 -114
rect 112 -322 146 -306
rect -100 -399 -84 -365
rect 84 -399 100 -365
rect -100 -507 -84 -473
rect 84 -507 100 -473
rect -146 -566 -112 -550
rect -146 -758 -112 -742
rect 112 -566 146 -550
rect 112 -758 146 -742
rect -100 -835 -84 -801
rect 84 -835 100 -801
rect -100 -943 -84 -909
rect 84 -943 100 -909
rect -146 -1002 -112 -986
rect -146 -1194 -112 -1178
rect 112 -1002 146 -986
rect 112 -1194 146 -1178
rect -100 -1271 -84 -1237
rect 84 -1271 100 -1237
rect -100 -1379 -84 -1345
rect 84 -1379 100 -1345
rect -146 -1438 -112 -1422
rect -146 -1630 -112 -1614
rect 112 -1438 146 -1422
rect 112 -1630 146 -1614
rect -100 -1707 -84 -1673
rect 84 -1707 100 -1673
rect -260 -1775 -226 -1713
rect 226 -1775 260 -1713
rect -260 -1809 -164 -1775
rect 164 -1809 260 -1775
<< viali >>
rect -84 1673 84 1707
rect -146 1438 -112 1614
rect 112 1438 146 1614
rect -84 1345 84 1379
rect -84 1237 84 1271
rect -146 1002 -112 1178
rect 112 1002 146 1178
rect -84 909 84 943
rect -84 801 84 835
rect -146 566 -112 742
rect 112 566 146 742
rect -84 473 84 507
rect -84 365 84 399
rect -146 130 -112 306
rect 112 130 146 306
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -306 -112 -130
rect 112 -306 146 -130
rect -84 -399 84 -365
rect -84 -507 84 -473
rect -146 -742 -112 -566
rect 112 -742 146 -566
rect -84 -835 84 -801
rect -84 -943 84 -909
rect -146 -1178 -112 -1002
rect 112 -1178 146 -1002
rect -84 -1271 84 -1237
rect -84 -1379 84 -1345
rect -146 -1614 -112 -1438
rect 112 -1614 146 -1438
rect -84 -1707 84 -1673
<< metal1 >>
rect -96 1707 96 1713
rect -96 1673 -84 1707
rect 84 1673 96 1707
rect -96 1667 96 1673
rect -152 1614 -106 1626
rect -152 1438 -146 1614
rect -112 1438 -106 1614
rect -152 1426 -106 1438
rect 106 1614 152 1626
rect 106 1438 112 1614
rect 146 1438 152 1614
rect 106 1426 152 1438
rect -96 1379 96 1385
rect -96 1345 -84 1379
rect 84 1345 96 1379
rect -96 1339 96 1345
rect -96 1271 96 1277
rect -96 1237 -84 1271
rect 84 1237 96 1271
rect -96 1231 96 1237
rect -152 1178 -106 1190
rect -152 1002 -146 1178
rect -112 1002 -106 1178
rect -152 990 -106 1002
rect 106 1178 152 1190
rect 106 1002 112 1178
rect 146 1002 152 1178
rect 106 990 152 1002
rect -96 943 96 949
rect -96 909 -84 943
rect 84 909 96 943
rect -96 903 96 909
rect -96 835 96 841
rect -96 801 -84 835
rect 84 801 96 835
rect -96 795 96 801
rect -152 742 -106 754
rect -152 566 -146 742
rect -112 566 -106 742
rect -152 554 -106 566
rect 106 742 152 754
rect 106 566 112 742
rect 146 566 152 742
rect 106 554 152 566
rect -96 507 96 513
rect -96 473 -84 507
rect 84 473 96 507
rect -96 467 96 473
rect -96 399 96 405
rect -96 365 -84 399
rect 84 365 96 399
rect -96 359 96 365
rect -152 306 -106 318
rect -152 130 -146 306
rect -112 130 -106 306
rect -152 118 -106 130
rect 106 306 152 318
rect 106 130 112 306
rect 146 130 152 306
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -306 -146 -130
rect -112 -306 -106 -130
rect -152 -318 -106 -306
rect 106 -130 152 -118
rect 106 -306 112 -130
rect 146 -306 152 -130
rect 106 -318 152 -306
rect -96 -365 96 -359
rect -96 -399 -84 -365
rect 84 -399 96 -365
rect -96 -405 96 -399
rect -96 -473 96 -467
rect -96 -507 -84 -473
rect 84 -507 96 -473
rect -96 -513 96 -507
rect -152 -566 -106 -554
rect -152 -742 -146 -566
rect -112 -742 -106 -566
rect -152 -754 -106 -742
rect 106 -566 152 -554
rect 106 -742 112 -566
rect 146 -742 152 -566
rect 106 -754 152 -742
rect -96 -801 96 -795
rect -96 -835 -84 -801
rect 84 -835 96 -801
rect -96 -841 96 -835
rect -96 -909 96 -903
rect -96 -943 -84 -909
rect 84 -943 96 -909
rect -96 -949 96 -943
rect -152 -1002 -106 -990
rect -152 -1178 -146 -1002
rect -112 -1178 -106 -1002
rect -152 -1190 -106 -1178
rect 106 -1002 152 -990
rect 106 -1178 112 -1002
rect 146 -1178 152 -1002
rect 106 -1190 152 -1178
rect -96 -1237 96 -1231
rect -96 -1271 -84 -1237
rect 84 -1271 96 -1237
rect -96 -1277 96 -1271
rect -96 -1345 96 -1339
rect -96 -1379 -84 -1345
rect 84 -1379 96 -1345
rect -96 -1385 96 -1379
rect -152 -1438 -106 -1426
rect -152 -1614 -146 -1438
rect -112 -1614 -106 -1438
rect -152 -1626 -106 -1614
rect 106 -1438 152 -1426
rect 106 -1614 112 -1438
rect 146 -1614 152 -1438
rect 106 -1626 152 -1614
rect -96 -1673 96 -1667
rect -96 -1707 -84 -1673
rect 84 -1707 96 -1673
rect -96 -1713 96 -1707
<< properties >>
string FIXED_BBOX -243 -1792 243 1792
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
