magic
tech sky130A
magscale 1 2
timestamp 1769859645
<< nwell >>
rect 1000 -600 2200 3200
<< viali >>
rect 1040 -3200 1380 -3140
rect 1640 -3200 1980 -3140
<< metal1 >>
rect 1000 3000 1800 3600
rect 1240 2900 1800 3000
rect 800 2800 1100 2900
rect 800 2600 1200 2800
rect 1000 1200 1400 2400
rect 1700 1200 1800 2900
rect 700 660 1340 720
rect 1880 700 2340 720
rect 1880 660 2480 700
rect 700 200 860 660
rect 1220 600 1300 620
rect 600 0 860 200
rect 700 -420 860 0
rect 900 560 1180 580
rect 900 -260 920 560
rect 1160 -260 1180 560
rect 900 -280 1180 -260
rect 1220 -360 1240 600
rect 1820 600 1900 620
rect 1360 520 1780 580
rect 1360 -260 1460 520
rect 1680 -260 1780 520
rect 1360 -360 1780 -260
rect 1820 -340 1840 600
rect 1960 520 2180 540
rect 1960 -220 1980 520
rect 2160 -220 2180 520
rect 1960 -240 2180 -220
rect 2260 200 2480 660
rect 2260 0 2600 200
rect 1820 -360 1900 -340
rect 1220 -380 1300 -360
rect 2260 -420 2480 0
rect 700 -480 1260 -420
rect 1780 -480 2480 -420
rect 2400 -620 2600 -600
rect 2400 -780 2420 -620
rect 2580 -780 2600 -620
rect 2400 -800 2600 -780
rect 900 -2760 1160 -1100
rect 900 -3120 1000 -2760
rect 1240 -3020 1320 -2400
rect 1860 -2880 2100 -1200
rect 1180 -3080 1860 -3020
rect 2000 -3120 2100 -2880
rect 900 -3140 2100 -3120
rect 900 -3200 1040 -3140
rect 1380 -3200 1640 -3140
rect 1980 -3200 2100 -3140
rect 600 -3400 2100 -3200
<< via1 >>
rect 920 -260 1160 560
rect 1240 -360 1300 600
rect 1460 -260 1680 520
rect 1840 -340 1900 600
rect 1980 -220 2160 520
rect 2420 -780 2580 -620
<< metal2 >>
rect 1000 1200 1400 2400
rect 1220 600 1300 620
rect 900 560 1180 580
rect 900 -260 920 560
rect 1160 -260 1180 560
rect 900 -280 1180 -260
rect 1220 -360 1240 600
rect 1820 600 1900 620
rect 1440 520 1700 540
rect 1440 -260 1460 520
rect 1680 -260 1700 520
rect 1440 -280 1700 -260
rect 1820 -340 1840 600
rect 1960 520 2180 540
rect 1960 -220 1980 520
rect 2160 -220 2180 520
rect 1960 -240 2180 -220
rect 1820 -360 1900 -340
rect 1220 -380 1300 -360
rect 1600 -620 2600 -600
rect 1600 -780 2420 -620
rect 2580 -780 2600 -620
rect 1600 -800 2600 -780
<< via2 >>
rect 920 -260 1160 560
rect 1460 -260 1680 520
rect 1980 -220 2160 520
<< metal3 >>
rect 1000 580 1400 2400
rect 900 560 1400 580
rect 900 -260 920 560
rect 1160 540 1720 560
rect 1160 520 2180 540
rect 1160 -260 1460 520
rect 1680 -220 1980 520
rect 2160 -220 2180 520
rect 1680 -260 2180 -220
rect 900 -280 1720 -260
use sky130_fd_pr__nfet_01v8_A5WNKR  sky130_fd_pr__nfet_01v8_A5WNKR_0
timestamp 1768764364
transform 1 0 1811 0 1 -2021
box -211 -1179 211 1179
use sky130_fd_pr__pfet_01v8_MGEV6J  sky130_fd_pr__pfet_01v8_MGEV6J_0
timestamp 1768764364
transform 1 0 1863 0 1 119
box -263 -719 263 719
use sky130_fd_pr__pfet_01v8_SB2EVP  XM1
timestamp 1769859645
transform 1 0 1496 0 1 1984
box -576 -4184 404 1256
use sky130_fd_pr__nfet_01v8_A5WNKR  XM2
timestamp 1768764364
transform 1 0 1211 0 1 -2021
box -211 -1179 211 1179
use sky130_fd_pr__pfet_01v8_MGEV6J  XM4
timestamp 1768764364
transform 1 0 1263 0 1 119
box -263 -719 263 719
<< labels >>
flabel metal1 600 -3400 800 -3200 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 1000 3400 1200 3600 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 800 2600 1000 2800 0 FreeSans 256 0 0 0 PBIAS
port 5 nsew
flabel metal1 600 0 800 200 0 FreeSans 256 0 0 0 AMP_P
port 3 nsew
flabel metal1 2400 0 2600 200 0 FreeSans 256 0 0 0 AMP_N
port 4 nsew
flabel metal1 2400 -800 2600 -600 0 FreeSans 256 0 0 0 AMP_OUT
port 2 nsew
<< end >>
