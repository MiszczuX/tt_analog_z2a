magic
tech sky130A
magscale 1 2
timestamp 1769859645
<< error_p >>
rect -476 396 -467 405
rect -125 396 -116 405
rect -485 391 -107 396
rect -485 387 -471 391
rect -476 -755 -471 387
rect -485 -759 -471 -755
rect -121 387 -107 391
rect -121 -755 -116 387
rect 278 -324 284 976
rect -121 -759 -107 -755
rect -485 -764 -107 -759
rect -476 -773 -467 -764
rect -125 -773 -116 -764
<< nwell >>
rect -296 -984 296 984
<< pmos >>
rect -100 -836 100 764
<< pdiff >>
rect -158 752 -100 764
rect -158 -824 -146 752
rect -112 -824 -100 752
rect -158 -836 -100 -824
rect 100 752 158 764
rect 100 -824 112 752
rect 146 -824 158 752
rect 100 -836 158 -824
<< pdiffc >>
rect -146 -824 -112 752
rect 112 -824 146 752
<< nsubdiff >>
rect -260 914 -164 948
rect 164 914 260 948
rect -260 851 -226 914
rect 226 851 260 914
rect -260 -914 -226 -851
rect 226 -914 260 -851
rect -260 -948 -164 -914
rect 164 -948 260 -914
<< nsubdiffcont >>
rect -164 914 164 948
rect -260 -851 -226 851
rect 226 -851 260 851
rect -164 -948 164 -914
<< poly >>
rect -100 845 100 861
rect -100 811 -84 845
rect 84 811 100 845
rect -100 764 100 811
rect -100 -862 100 -836
<< polycont >>
rect -84 811 84 845
<< locali >>
rect -260 914 -164 948
rect 164 914 204 948
rect -260 851 -226 914
rect -100 811 -84 845
rect 84 811 100 845
rect -146 752 -112 768
rect -146 -840 -112 -824
rect 112 752 146 768
rect 112 -840 146 -824
rect -260 -914 -226 -851
rect 226 -914 260 -851
rect -260 -948 -164 -914
rect 164 -948 260 -914
<< viali >>
rect 204 851 284 976
rect -84 811 84 845
rect -146 -824 -112 752
rect 112 -824 146 752
rect 204 -324 226 851
rect 226 -324 260 851
rect 260 -324 284 851
<< metal1 >>
rect 164 976 284 1256
rect -576 851 4 856
rect -576 845 96 851
rect -576 811 -84 845
rect 84 811 96 845
rect -576 805 96 811
rect -576 796 4 805
rect 164 796 204 976
rect 124 764 204 796
rect -152 752 -106 764
rect -152 396 -146 752
rect -152 -824 -146 -764
rect -112 -824 -106 752
rect -152 -836 -106 -824
rect 106 752 204 764
rect 106 -824 112 752
rect 146 -324 204 752
rect 146 -784 284 -324
rect 146 -824 152 -784
rect 106 -836 152 -824
rect -256 -3104 -96 -3084
rect -256 -4144 -196 -3104
rect -116 -4144 -96 -3104
rect -256 -4184 -96 -4144
rect 104 -3124 304 -3084
rect 104 -4164 144 -3124
rect 224 -4164 304 -3124
rect 104 -4184 304 -4164
<< via1 >>
rect -476 -764 -146 396
rect -146 -764 -116 396
rect -196 -4144 -116 -3104
rect 144 -4164 224 -3124
<< metal2 >>
rect -296 -2384 -196 -2284
rect 304 -2384 404 -2284
rect -296 -2484 -96 -2384
rect -196 -3084 -96 -2484
rect -236 -3104 -96 -3084
rect -236 -4144 -196 -3104
rect -116 -4144 -96 -3104
rect -236 -4184 -96 -4144
rect 104 -2484 404 -2384
rect 104 -3084 204 -2484
rect 104 -3124 244 -3084
rect 104 -4164 144 -3124
rect 224 -4164 244 -3124
rect 104 -4184 244 -4164
<< via2 >>
rect -476 -764 -116 396
<< properties >>
string FIXED_BBOX -243 -931 243 931
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
