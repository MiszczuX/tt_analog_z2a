magic
tech sky130A
magscale 1 2
timestamp 1765032183
<< metal1 >>
rect 25704 3086 25710 3286
rect 25910 3086 27330 3286
rect 30600 2516 30800 2522
rect 26480 2316 26486 2516
rect 26686 2316 27330 2516
rect 30600 2310 30800 2316
rect 25902 1626 25908 1826
rect 26108 1626 27356 1826
<< via1 >>
rect 25710 3086 25910 3286
rect 26486 2316 26686 2516
rect 30600 2316 30800 2516
rect 25908 1626 26108 1826
<< metal2 >>
rect 25710 3286 25910 3292
rect 25701 3086 25710 3286
rect 25910 3086 25919 3286
rect 25710 3080 25910 3086
rect 26486 2516 26686 2525
rect 30600 2516 30800 2525
rect 30594 2316 30600 2516
rect 30800 2316 30806 2516
rect 26486 2307 26686 2316
rect 30600 2307 30800 2316
rect 25908 1826 26108 1832
rect 25899 1626 25908 1826
rect 26108 1626 26117 1826
rect 25908 1620 26108 1626
<< via2 >>
rect 25710 3086 25910 3286
rect 26486 2316 26686 2516
rect 30600 2316 30800 2516
rect 25908 1626 26108 1826
<< metal3 >>
rect 324 3286 524 3292
rect 25705 3286 25915 3291
rect 524 3086 25710 3286
rect 25910 3086 25915 3286
rect 324 3080 524 3086
rect 25705 3081 25915 3086
rect 26481 2516 26691 2521
rect 26481 2511 26486 2516
rect 26686 2511 26691 2516
rect 26481 2305 26691 2311
rect 30595 2516 30805 2521
rect 30595 2511 30600 2516
rect 30800 2511 30805 2516
rect 30595 2305 30805 2311
rect 25897 1621 25903 1831
rect 26103 1826 26113 1831
rect 26108 1626 26113 1826
rect 26103 1621 26113 1626
<< via3 >>
rect 324 3086 524 3286
rect 26481 2316 26486 2511
rect 26486 2316 26686 2511
rect 26686 2316 26691 2511
rect 26481 2311 26691 2316
rect 30595 2316 30600 2511
rect 30600 2316 30800 2511
rect 30800 2316 30805 2511
rect 30595 2311 30805 2316
rect 25903 1826 26103 1831
rect 25903 1626 25908 1826
rect 25908 1626 26103 1826
rect 25903 1621 26103 1626
<< metal4 >>
rect 200 3286 600 44152
rect 200 3086 324 3286
rect 524 3086 600 3286
rect 200 1000 600 3086
rect 800 42376 1200 44152
rect 6134 42376 6194 45152
rect 6686 42376 6746 45152
rect 7238 42376 7298 45152
rect 7790 42376 7850 45152
rect 8342 42376 8402 45152
rect 8894 42376 8954 45152
rect 9446 42376 9506 45152
rect 9998 42376 10058 45152
rect 10550 42376 10610 45152
rect 11102 42376 11162 45152
rect 11654 42376 11714 45152
rect 12206 42376 12266 45152
rect 12758 42376 12818 45152
rect 13310 42376 13370 45152
rect 13862 42376 13922 45152
rect 14414 42376 14474 45152
rect 14966 42376 15026 45152
rect 15518 42376 15578 45152
rect 16070 42376 16130 45152
rect 16622 42376 16682 45152
rect 17174 42376 17234 45152
rect 17726 42376 17786 45152
rect 18278 42376 18338 45152
rect 18830 45014 18890 45152
rect 18826 42376 18894 45014
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 800 42308 18894 42376
rect 800 1826 1200 42308
rect 26480 2511 26692 2512
rect 26480 2311 26481 2511
rect 26691 2311 26692 2511
rect 26480 2310 26692 2311
rect 30594 2511 30806 2512
rect 30594 2311 30595 2511
rect 30805 2311 30806 2511
rect 30594 2310 30806 2311
rect 25902 1831 26104 1832
rect 25902 1826 25903 1831
rect 800 1626 25903 1826
rect 800 1000 1200 1626
rect 25902 1621 25903 1626
rect 26103 1621 26104 1831
rect 25902 1620 26104 1621
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26486 48 26686 2310
rect 30600 1150 30800 2310
rect 30344 950 30800 1150
rect 30344 510 30544 950
rect 26498 0 26678 48
rect 30362 0 30542 510
use double_inverter  double_inverter_0
timestamp 1764265104
transform 1 0 25970 0 1 3086
box 1160 -1520 4830 250
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
