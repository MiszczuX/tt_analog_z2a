magic
tech sky130A
magscale 1 2
timestamp 1764261594
<< error_p >>
rect -365 181 -307 187
rect -173 181 -115 187
rect 19 181 77 187
rect 211 181 269 187
rect 403 181 461 187
rect -365 147 -353 181
rect -173 147 -161 181
rect 19 147 31 181
rect 211 147 223 181
rect 403 147 415 181
rect -365 141 -307 147
rect -173 141 -115 147
rect 19 141 77 147
rect 211 141 269 147
rect 403 141 461 147
rect -461 -147 -403 -141
rect -269 -147 -211 -141
rect -77 -147 -19 -141
rect 115 -147 173 -141
rect 307 -147 365 -141
rect -461 -181 -449 -147
rect -269 -181 -257 -147
rect -77 -181 -65 -147
rect 115 -181 127 -147
rect 307 -181 319 -147
rect -461 -187 -403 -181
rect -269 -187 -211 -181
rect -77 -187 -19 -181
rect 115 -187 173 -181
rect 307 -187 365 -181
<< nwell >>
rect -647 -319 647 319
<< pmos >>
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
<< pdiff >>
rect -509 88 -447 100
rect -509 -88 -497 88
rect -463 -88 -447 88
rect -509 -100 -447 -88
rect -417 88 -351 100
rect -417 -88 -401 88
rect -367 -88 -351 88
rect -417 -100 -351 -88
rect -321 88 -255 100
rect -321 -88 -305 88
rect -271 -88 -255 88
rect -321 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 321 100
rect 255 -88 271 88
rect 305 -88 321 88
rect 255 -100 321 -88
rect 351 88 417 100
rect 351 -88 367 88
rect 401 -88 417 88
rect 351 -100 417 -88
rect 447 88 509 100
rect 447 -88 463 88
rect 497 -88 509 88
rect 447 -100 509 -88
<< pdiffc >>
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
<< nsubdiff >>
rect -611 249 -515 283
rect 515 249 611 283
rect -611 187 -577 249
rect 577 187 611 249
rect -611 -249 -577 -187
rect 577 -249 611 -187
rect -611 -283 -515 -249
rect 515 -283 611 -249
<< nsubdiffcont >>
rect -515 249 515 283
rect -611 -187 -577 187
rect 577 -187 611 187
rect -515 -283 515 -249
<< poly >>
rect -369 181 -303 197
rect -369 147 -353 181
rect -319 147 -303 181
rect -369 131 -303 147
rect -177 181 -111 197
rect -177 147 -161 181
rect -127 147 -111 181
rect -177 131 -111 147
rect 15 181 81 197
rect 15 147 31 181
rect 65 147 81 181
rect 15 131 81 147
rect 207 181 273 197
rect 207 147 223 181
rect 257 147 273 181
rect 207 131 273 147
rect 399 181 465 197
rect 399 147 415 181
rect 449 147 465 181
rect 399 131 465 147
rect -447 100 -417 126
rect -351 100 -321 131
rect -255 100 -225 126
rect -159 100 -129 131
rect -63 100 -33 126
rect 33 100 63 131
rect 129 100 159 126
rect 225 100 255 131
rect 321 100 351 126
rect 417 100 447 131
rect -447 -131 -417 -100
rect -351 -126 -321 -100
rect -255 -131 -225 -100
rect -159 -126 -129 -100
rect -63 -131 -33 -100
rect 33 -126 63 -100
rect 129 -131 159 -100
rect 225 -126 255 -100
rect 321 -131 351 -100
rect 417 -126 447 -100
rect -465 -147 -399 -131
rect -465 -181 -449 -147
rect -415 -181 -399 -147
rect -465 -197 -399 -181
rect -273 -147 -207 -131
rect -273 -181 -257 -147
rect -223 -181 -207 -147
rect -273 -197 -207 -181
rect -81 -147 -15 -131
rect -81 -181 -65 -147
rect -31 -181 -15 -147
rect -81 -197 -15 -181
rect 111 -147 177 -131
rect 111 -181 127 -147
rect 161 -181 177 -147
rect 111 -197 177 -181
rect 303 -147 369 -131
rect 303 -181 319 -147
rect 353 -181 369 -147
rect 303 -197 369 -181
<< polycont >>
rect -353 147 -319 181
rect -161 147 -127 181
rect 31 147 65 181
rect 223 147 257 181
rect 415 147 449 181
rect -449 -181 -415 -147
rect -257 -181 -223 -147
rect -65 -181 -31 -147
rect 127 -181 161 -147
rect 319 -181 353 -147
<< locali >>
rect -611 249 -515 283
rect 515 249 611 283
rect -611 187 -577 249
rect 577 187 611 249
rect -369 147 -353 181
rect -319 147 -303 181
rect -177 147 -161 181
rect -127 147 -111 181
rect 15 147 31 181
rect 65 147 81 181
rect 207 147 223 181
rect 257 147 273 181
rect 399 147 415 181
rect 449 147 465 181
rect -497 88 -463 104
rect -497 -104 -463 -88
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect 463 88 497 104
rect 463 -104 497 -88
rect -465 -181 -449 -147
rect -415 -181 -399 -147
rect -273 -181 -257 -147
rect -223 -181 -207 -147
rect -81 -181 -65 -147
rect -31 -181 -15 -147
rect 111 -181 127 -147
rect 161 -181 177 -147
rect 303 -181 319 -147
rect 353 -181 369 -147
rect -611 -249 -577 -187
rect 577 -249 611 -187
rect -611 -283 -515 -249
rect 515 -283 611 -249
<< viali >>
rect -353 147 -319 181
rect -161 147 -127 181
rect 31 147 65 181
rect 223 147 257 181
rect 415 147 449 181
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect -449 -181 -415 -147
rect -257 -181 -223 -147
rect -65 -181 -31 -147
rect 127 -181 161 -147
rect 319 -181 353 -147
<< metal1 >>
rect -365 181 -307 187
rect -365 147 -353 181
rect -319 147 -307 181
rect -365 141 -307 147
rect -173 181 -115 187
rect -173 147 -161 181
rect -127 147 -115 181
rect -173 141 -115 147
rect 19 181 77 187
rect 19 147 31 181
rect 65 147 77 181
rect 19 141 77 147
rect 211 181 269 187
rect 211 147 223 181
rect 257 147 269 181
rect 211 141 269 147
rect 403 181 461 187
rect 403 147 415 181
rect 449 147 461 181
rect 403 141 461 147
rect -503 88 -457 100
rect -503 -88 -497 88
rect -463 -88 -457 88
rect -503 -100 -457 -88
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
rect 457 88 503 100
rect 457 -88 463 88
rect 497 -88 503 88
rect 457 -100 503 -88
rect -461 -147 -403 -141
rect -461 -181 -449 -147
rect -415 -181 -403 -147
rect -461 -187 -403 -181
rect -269 -147 -211 -141
rect -269 -181 -257 -147
rect -223 -181 -211 -147
rect -269 -187 -211 -181
rect -77 -147 -19 -141
rect -77 -181 -65 -147
rect -31 -181 -19 -147
rect -77 -187 -19 -181
rect 115 -147 173 -141
rect 115 -181 127 -147
rect 161 -181 173 -147
rect 115 -187 173 -181
rect 307 -147 365 -141
rect 307 -181 319 -147
rect 353 -181 365 -147
rect 307 -187 365 -181
<< properties >>
string FIXED_BBOX -594 -266 594 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
