magic
tech sky130A
timestamp 1769869012
<< metal1 >>
rect 480000 561800 480700 562000
rect 490200 561900 492000 562000
rect 480000 560200 480200 561800
rect 491300 561650 491600 561700
rect 490400 561400 491000 561500
rect 491300 561250 491350 561650
rect 491550 561250 491600 561650
rect 491300 561200 491600 561250
rect 492500 561100 492900 562000
rect 494800 561870 495000 561900
rect 494800 561220 494820 561870
rect 494980 561220 495000 561870
rect 494800 561200 495000 561220
rect 490200 561000 490450 561100
rect 487400 560950 490450 561000
rect 490950 561000 491100 561100
rect 490950 560950 491300 561000
rect 487400 560900 491300 560950
rect 480000 560000 480700 560200
rect 480000 559600 482300 560000
rect 488100 559800 488400 560900
rect 492900 560650 493200 560700
rect 492900 560350 492950 560650
rect 493150 560350 493200 560650
rect 492900 560300 493200 560350
rect 480000 558800 482700 559600
rect 484600 559500 488400 559800
rect 494800 559700 495000 560200
rect 484600 558800 484800 559500
rect 485100 558900 488800 559100
rect 492600 559000 494800 559100
rect 492800 558900 494800 559000
rect 480000 557900 482300 558800
rect 484300 558700 484400 558800
rect 485100 558700 485300 558900
rect 484300 558500 485300 558700
rect 488500 558500 488800 558900
rect 494500 558000 494800 558900
rect 491300 557700 494800 558000
rect 492400 556300 493800 556600
rect 493400 556200 493800 556300
rect 493400 549600 493700 556200
rect 493500 549400 493700 549600
rect 479700 548200 480200 548300
rect 479700 548100 480000 548200
rect 480050 548100 480200 548200
rect 482500 546100 482750 546500
rect 483150 543750 483600 543800
rect 483150 543650 483200 543750
rect 483550 543650 483600 543750
rect 483150 543600 483600 543650
rect 493000 543600 493700 543700
rect 482300 543530 483100 543550
rect 480000 543450 482200 543500
rect 480000 543150 480200 543450
rect 480000 542150 480050 543150
rect 480150 542150 480200 543150
rect 480000 542100 480200 542150
rect 480300 543350 482000 543400
rect 480300 543150 480500 543350
rect 480300 542150 480350 543150
rect 480450 542150 480500 543150
rect 480300 542100 480500 542150
rect 480600 543250 481800 543300
rect 480600 543150 480800 543250
rect 480600 542150 480650 543150
rect 480750 542150 480800 543150
rect 480600 542100 480800 542150
rect 480900 543150 481600 543200
rect 480900 542150 480950 543150
rect 481050 543050 481600 543150
rect 481700 543050 481800 543250
rect 481900 543100 482000 543350
rect 482100 543100 482200 543450
rect 482300 543420 482580 543530
rect 483070 543420 483100 543530
rect 482300 543400 483100 543420
rect 482300 543100 482400 543400
rect 482500 543300 484250 543350
rect 482500 543100 482600 543300
rect 482700 543200 483950 543250
rect 482700 543100 482800 543200
rect 482900 543100 483650 543150
rect 481050 542150 481100 543050
rect 482500 542682 482600 543000
rect 483150 542900 483350 542950
rect 483150 542400 483200 542900
rect 480900 542100 481100 542150
rect 481200 542100 481350 542400
rect 483050 542200 483200 542400
rect 483300 542200 483350 542900
rect 483050 542150 483350 542200
rect 483450 542200 483500 543100
rect 483600 542200 483650 543100
rect 483450 542150 483650 542200
rect 483750 543100 483950 543200
rect 483750 542200 483800 543100
rect 483900 542200 483950 543100
rect 483750 542150 483950 542200
rect 484050 543200 484250 543300
rect 484050 542200 484100 543200
rect 484200 542200 484250 543200
rect 493000 543100 493200 543600
rect 493600 543100 493700 543600
rect 493000 543000 493700 543100
rect 493600 542800 493700 543000
rect 494500 542600 494800 557700
rect 484050 542150 484250 542200
rect 481250 542000 484900 542100
rect 491400 541800 492100 542500
rect 492200 542000 494800 542600
<< via1 >>
rect 491350 561250 491550 561650
rect 494820 561220 494980 561870
rect 490450 560950 490950 561100
rect 492950 560350 493150 560650
rect 483200 543650 483550 543750
rect 480050 542150 480150 543150
rect 480350 542150 480450 543150
rect 480650 542150 480750 543150
rect 480950 542150 481050 543150
rect 482580 543420 483070 543530
rect 483200 542200 483300 542900
rect 483500 542200 483600 543100
rect 483800 542200 483900 543100
rect 484100 542200 484200 543200
rect 493200 543100 493600 543600
<< metal2 >>
rect 494800 561870 495000 561900
rect 491300 561650 491600 561700
rect 480000 561300 480500 561600
rect 480000 558700 480200 561300
rect 491300 561250 491350 561650
rect 491550 561250 491600 561650
rect 491300 561200 491600 561250
rect 494800 561220 494820 561870
rect 494980 561220 495000 561870
rect 494800 561200 495000 561220
rect 490400 560950 490450 561100
rect 490950 560950 493200 561100
rect 490400 560900 493200 560950
rect 487800 560400 492700 560700
rect 492500 559300 492700 560400
rect 492900 560650 493200 560900
rect 492900 560350 492950 560650
rect 493150 560350 493200 560650
rect 492900 560300 493200 560350
rect 480000 558500 485500 558700
rect 492500 558400 492800 559300
rect 493000 556900 493200 560300
rect 493300 558700 493400 560100
rect 494800 559700 495000 560200
rect 493800 558800 494300 558900
rect 493300 558600 493600 558700
rect 493300 558300 493400 558600
rect 493500 558300 493600 558600
rect 493800 558600 493900 558800
rect 494200 558600 494300 558800
rect 493800 558500 494300 558600
rect 493300 558200 493600 558300
rect 492000 555700 493200 556900
rect 493900 556200 494200 558500
rect 493900 550700 494400 550800
rect 493900 550400 494000 550700
rect 494300 550400 494400 550700
rect 493900 550300 494400 550400
rect 482500 546100 482750 546500
rect 479800 544100 480500 544300
rect 480000 543150 480200 543200
rect 480000 542150 480050 543150
rect 480150 542150 480200 543150
rect 480000 542100 480200 542150
rect 480300 543150 480500 544100
rect 482300 543550 482400 544000
rect 483150 543750 483600 543800
rect 483150 543650 483200 543750
rect 483550 543650 483600 543750
rect 483150 543600 483600 543650
rect 492200 543600 493700 543700
rect 482300 543530 483100 543550
rect 482300 543420 482580 543530
rect 483070 543420 483100 543530
rect 482300 543400 483100 543420
rect 480300 542150 480350 543150
rect 480450 542150 480500 543150
rect 480300 542100 480500 542150
rect 480600 543150 480800 543200
rect 480600 542150 480650 543150
rect 480750 542150 480800 543150
rect 480600 542100 480800 542150
rect 480900 543150 481100 543200
rect 480900 542150 480950 543150
rect 481050 542150 481100 543150
rect 483150 542900 483350 543600
rect 484050 543200 484250 543250
rect 483150 542200 483200 542900
rect 483300 542200 483350 542900
rect 483150 542150 483350 542200
rect 483450 543100 483650 543150
rect 483450 542200 483500 543100
rect 483600 542200 483650 543100
rect 483450 542150 483650 542200
rect 483750 543100 483950 543150
rect 483750 542200 483800 543100
rect 483900 542200 483950 543100
rect 483750 542150 483950 542200
rect 484050 542200 484100 543200
rect 484200 542200 484250 543200
rect 484050 542150 484250 542200
rect 492200 543100 493200 543600
rect 493600 543100 493700 543600
rect 492200 543000 493700 543100
rect 480900 542100 481100 542150
rect 492200 542000 493500 543000
<< via2 >>
rect 491350 561250 491550 561650
rect 494820 561220 494980 561870
rect 493400 558300 493500 558600
rect 493900 558600 494200 558800
rect 494000 550400 494300 550700
rect 480050 542150 480150 543150
rect 480650 542150 480750 543150
rect 480950 542150 481050 543150
rect 483500 542200 483600 543100
rect 483800 542200 483900 543100
rect 484100 542200 484200 543200
<< metal3 >>
rect 494800 561870 495000 561900
rect 494800 561800 494820 561870
rect 491300 561650 491600 561700
rect 491300 561250 491350 561650
rect 491550 561250 491600 561650
rect 491300 561200 491600 561250
rect 491400 560700 491600 561200
rect 487500 560400 491600 560700
rect 491700 561300 494820 561800
rect 487500 559400 487800 560400
rect 491700 560000 492000 561300
rect 494800 561220 494820 561300
rect 494980 561220 495000 561870
rect 494800 561200 495000 561220
rect 486500 559100 487800 559400
rect 489500 559600 492000 560000
rect 486500 558500 486800 559100
rect 487500 557500 487800 558700
rect 489500 558300 489800 559600
rect 490500 558900 494300 559300
rect 490500 558600 490800 558900
rect 493800 558800 494300 558900
rect 491400 558000 491900 558700
rect 492800 558600 493600 558700
rect 492800 558300 493400 558600
rect 493500 558300 493600 558600
rect 493800 558600 493900 558800
rect 494200 558600 494300 558800
rect 493800 558500 494300 558600
rect 492800 558200 493600 558300
rect 494800 558000 495000 560200
rect 491400 557800 495000 558000
rect 487500 557300 493300 557500
rect 493000 550800 493300 557300
rect 493000 550700 494400 550800
rect 493000 550400 494000 550700
rect 494300 550400 494400 550700
rect 493000 550300 494400 550400
rect 483700 548200 484250 548650
rect 482500 546460 482750 546500
rect 482500 546140 482540 546460
rect 482720 546140 482750 546460
rect 482500 546100 482750 546140
rect 481200 543800 481300 546000
rect 483700 544550 483800 546000
rect 481200 543700 482500 543800
rect 480000 543150 480200 543200
rect 480000 542150 480050 543150
rect 480150 542150 480200 543150
rect 480000 542100 480200 542150
rect 480600 543150 480800 543200
rect 480600 542150 480650 543150
rect 480750 542150 480800 543150
rect 480600 542100 480800 542150
rect 480900 543150 481100 543200
rect 480900 542150 480950 543150
rect 481050 542150 481100 543150
rect 480900 542100 481100 542150
rect 482400 542100 482500 543700
rect 483700 543600 483950 544550
rect 483450 543350 483950 543600
rect 483450 543100 483650 543350
rect 484050 543200 484250 548200
rect 483450 542200 483500 543100
rect 483600 542200 483650 543100
rect 483450 542150 483650 542200
rect 483750 543100 483950 543150
rect 483750 542200 483800 543100
rect 483900 542200 483950 543100
rect 483750 542100 483950 542200
rect 484050 542200 484100 543200
rect 484200 542200 484250 543200
rect 484050 542150 484250 542200
rect 482400 542000 483950 542100
<< via3 >>
rect 482540 546140 482720 546460
rect 480050 542150 480150 543150
rect 480650 542150 480750 543150
rect 480950 542150 481050 543150
<< metal4 >>
rect 482300 546460 482750 546500
rect 482300 546140 482540 546460
rect 482720 546140 482750 546460
rect 482300 546100 482750 546140
rect 482300 545500 482500 546100
rect 482200 545300 482500 545500
rect 479700 543200 479800 544400
rect 480000 543400 480200 544400
rect 480300 543600 480500 544400
rect 480300 543500 481100 543600
rect 480000 543300 480800 543400
rect 479700 543150 480200 543200
rect 479700 542150 480050 543150
rect 480150 542150 480200 543150
rect 479700 542100 480200 542150
rect 480600 543150 480800 543300
rect 480600 542150 480650 543150
rect 480750 542150 480800 543150
rect 480600 542100 480800 542150
rect 480900 543150 481100 543500
rect 480900 542150 480950 543150
rect 481050 542150 481100 543150
rect 480900 542100 481100 542150
rect 482200 541800 482400 545300
use BG  BG_0
timestamp 1769856845
transform -1 0 483600 0 -1 541982
box 300 -1150 2400 -218
use BG  BG_1
timestamp 1769856845
transform 1 0 482300 0 1 559950
box 300 -1150 2400 -218
use inv_x1  inv_x1_0 ~/tt_analog_z2a_2/mag
timestamp 1769862601
transform 1 0 490900 0 1 561700
box 100 -700 500 200
use OSC3  OSC3_0 ~/tt_analog_z2a_2/mag
timestamp 1769852641
transform 0 1 494100 -1 0 556650
box 100 -500 4750 500
use OSC5  OSC5_0
timestamp 1769852641
transform 1 0 480400 0 -1 560500
box -100 -500 7500 500
use OSC5cap  OSC5cap_0
timestamp 1769636617
transform 0 1 494000 -1 0 550600
box 0 -800 7600 600
use OSC7  OSC7_0
timestamp 1769635987
transform 1 0 480200 0 1 561500
box 100 -500 10500 500
use T_FLIP_FLOP  T_FLIP_FLOP_0
timestamp 1769863106
transform 1 0 491600 0 1 561000
box 400 -2000 3400 1000
use VCMUX  VCMUX_0
timestamp 1769869012
transform 1 0 479400 0 1 547500
box -300 -5900 14100 11200
<< labels >>
rlabel metal1 480000 561900 480100 562000 1 VDD
port 4 n
rlabel metal1 493600 542800 493700 542900 1 VSS
port 2 n
rlabel metal1 492000 541800 492100 541900 1 VCMUXOUT
port 1 n
rlabel metal1 479900 548100 480000 548200 1 VCMUXIN
port 3 n
<< end >>
