magic
tech sky130A
magscale 1 2
timestamp 1770840455
<< pwell >>
rect 1000 -1900 5400 -500
<< viali >>
rect 5400 -1300 5440 -720
<< metal1 >>
rect 800 -1100 1300 -700
rect 1700 -1100 2200 -700
rect 2700 -1100 3300 -700
rect 3700 -1100 4300 -700
rect 4700 -1100 5300 -700
rect 5360 -720 5700 -700
rect 800 -1900 1000 -1100
rect 1200 -1700 1800 -1400
rect 1400 -2200 1600 -1700
rect 1900 -2200 2100 -1100
rect 2200 -1700 2800 -1300
rect 2400 -2200 2600 -1700
rect 2900 -2200 3100 -1100
rect 3200 -1700 3800 -1300
rect 3400 -2200 3600 -1700
rect 3900 -2200 4100 -1100
rect 4200 -1700 4800 -1300
rect 4400 -2200 4600 -1700
rect 4900 -2200 5100 -1100
rect 5360 -1300 5400 -720
rect 5440 -1300 5700 -720
rect 5200 -1700 5700 -1300
rect 5500 -1900 5700 -1700
use sky130_fd_pr__res_xhigh_po_0p69_87HR5C  XR0
timestamp 1770840455
transform 1 0 1235 0 1 -1218
box -235 -682 235 682
use sky130_fd_pr__res_xhigh_po_0p69_87HR5C  XR1
timestamp 1770840455
transform 1 0 1735 0 1 -1218
box -235 -682 235 682
use sky130_fd_pr__res_xhigh_po_0p69_87HR5C  XR2
timestamp 1770840455
transform 1 0 2235 0 1 -1218
box -235 -682 235 682
use sky130_fd_pr__res_xhigh_po_0p69_87HR5C  XR3
timestamp 1770840455
transform 1 0 2735 0 1 -1218
box -235 -682 235 682
use sky130_fd_pr__res_xhigh_po_0p69_87HR5C  XR4
timestamp 1770840455
transform 1 0 3235 0 1 -1218
box -235 -682 235 682
use sky130_fd_pr__res_xhigh_po_0p69_87HR5C  XR5
timestamp 1770840455
transform 1 0 3735 0 1 -1218
box -235 -682 235 682
use sky130_fd_pr__res_xhigh_po_0p69_87HR5C  XR6
timestamp 1770840455
transform 1 0 4235 0 1 -1218
box -235 -682 235 682
use sky130_fd_pr__res_xhigh_po_0p69_87HR5C  XR7
timestamp 1770840455
transform 1 0 4735 0 1 -1218
box -235 -682 235 682
use sky130_fd_pr__res_xhigh_po_0p69_87HR5C  XR8
timestamp 1770840455
transform 1 0 5235 0 1 -1218
box -235 -682 235 682
<< labels >>
flabel metal1 5500 -1900 5700 -1700 0 FreeSans 256 0 0 0 VSS
port 9 nsew
flabel metal1 4900 -2200 5100 -2000 0 FreeSans 256 0 0 0 vbg_0_2
port 7 nsew
flabel metal1 4400 -2200 4600 -2000 0 FreeSans 256 0 0 0 vbg_0_4
port 6 nsew
flabel metal1 3900 -2200 4100 -2000 0 FreeSans 256 0 0 0 vbg_0_6
port 5 nsew
flabel metal1 3400 -2200 3600 -2000 0 FreeSans 256 0 0 0 vbg_0_8
port 4 nsew
flabel metal1 2900 -2200 3100 -2000 0 FreeSans 256 0 0 0 vbg_1_0
port 3 nsew
flabel metal1 2400 -2200 2600 -2000 0 FreeSans 256 0 0 0 vbg_1_2
port 2 nsew
flabel metal1 1900 -2200 2100 -2000 0 FreeSans 256 0 0 0 vbg_1_4
port 1 nsew
flabel metal1 1400 -2200 1600 -2000 0 FreeSans 256 0 0 0 vbg_1_6
port 0 nsew
flabel metal1 800 -1900 1000 -1700 0 FreeSans 256 0 0 0 VDD
port 8 nsew
<< end >>
