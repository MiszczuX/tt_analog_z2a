** sch_path: /home/ttuser/tt_analog_z2a/xschem/PASSGATE.sch
.subckt PASSGATE VDD PASS_GATE_IN VSS PASS_GATE_EN PASS_GATE_OUT
*.PININFO PASS_GATE_IN:B PASS_GATE_EN:I VDD:B VSS:B PASS_GATE_OUT:B
XM1pass PASS_GATE_ZEN PASS_GATE_EN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=10 nf=1 m=1
XM0pass PASS_GATE_ZEN PASS_GATE_EN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 m=1
XM1 PASS_GATE_IN PASS_GATE_EN PASS_GATE_OUT VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 PASS_GATE_OUT PASS_GATE_ZEN PASS_GATE_IN VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends
.end
