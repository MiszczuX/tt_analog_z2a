magic
tech sky130A
magscale 1 2
timestamp 1768761543
<< error_p >>
rect -61 1018 -27 1024
rect -61 -946 -55 1018
rect -33 -946 -27 1018
rect -61 -952 -27 -946
rect -29 -1011 29 -1005
rect -29 -1045 -17 -1011
rect -29 -1051 29 -1045
<< nwell >>
rect -211 -1184 211 1184
<< pmos >>
rect -15 -964 15 1036
<< pdiff >>
rect -73 1024 -15 1036
rect -73 -952 -61 1024
rect -27 -952 -15 1024
rect -73 -964 -15 -952
rect 15 1024 73 1036
rect 15 -952 27 1024
rect 61 -952 73 1024
rect 15 -964 73 -952
<< pdiffc >>
rect -61 -952 -27 1024
rect 27 -952 61 1024
<< nsubdiff >>
rect -175 1114 -79 1148
rect 79 1114 175 1148
rect -175 1051 -141 1114
rect 141 1051 175 1114
rect -175 -1114 -141 -1051
rect 141 -1114 175 -1051
rect -175 -1148 -79 -1114
rect 79 -1148 175 -1114
<< nsubdiffcont >>
rect -79 1114 79 1148
rect -175 -1051 -141 1051
rect 141 -1051 175 1051
rect -79 -1148 79 -1114
<< poly >>
rect -15 1036 15 1062
rect -15 -995 15 -964
rect -33 -1011 33 -995
rect -33 -1045 -17 -1011
rect 17 -1045 33 -1011
rect -33 -1061 33 -1045
<< polycont >>
rect -17 -1045 17 -1011
<< locali >>
rect -175 1114 -79 1148
rect 79 1114 175 1148
rect -175 1051 -141 1114
rect 141 1051 175 1114
rect -61 1024 -27 1040
rect -61 -968 -27 -952
rect 27 1024 61 1040
rect 27 -968 61 -952
rect -33 -1045 -17 -1011
rect 17 -1045 33 -1011
rect -175 -1114 -141 -1051
rect 141 -1114 175 -1051
rect -175 -1148 -79 -1114
rect 79 -1148 175 -1114
<< viali >>
rect -61 -952 -27 1024
rect 27 -952 61 1024
rect -17 -1045 17 -1011
<< metal1 >>
rect 21 1024 67 1036
rect 21 -952 27 1024
rect 61 -952 67 1024
rect 21 -964 67 -952
rect -29 -1011 29 -1005
rect -29 -1045 -17 -1011
rect 17 -1045 29 -1011
rect -29 -1051 29 -1045
<< properties >>
string FIXED_BBOX -158 -1131 158 1131
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
