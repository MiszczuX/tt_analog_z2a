magic
tech sky130A
magscale 1 2
timestamp 1770560933
<< nwell >>
rect 600 400 1100 1600
<< viali >>
rect 680 1500 960 1560
rect 660 900 960 1060
rect 660 -400 960 -240
rect 660 -900 960 -840
<< metal1 >>
rect -200 1600 1000 1800
rect 600 1560 1000 1600
rect 600 1500 680 1560
rect 960 1500 1000 1560
rect 600 1480 1000 1500
rect 600 1400 780 1420
rect 600 1260 620 1400
rect 760 1260 780 1400
rect 600 1240 780 1260
rect 840 1220 1000 1480
rect 0 1180 560 1200
rect 0 1120 880 1180
rect 0 1100 560 1120
rect 0 200 100 1100
rect 640 1060 980 1080
rect 640 900 660 1060
rect 960 900 980 1060
rect 640 880 980 900
rect 600 800 780 820
rect 600 640 620 800
rect 760 640 780 800
rect 600 620 780 640
rect 840 620 980 880
rect 200 580 540 600
rect 200 420 220 580
rect 520 520 880 580
rect 520 420 540 520
rect 200 400 540 420
rect 1000 380 1200 400
rect 1000 220 1020 380
rect 1180 220 1200 380
rect 1000 200 1200 220
rect -200 140 400 200
rect -200 80 880 140
rect -200 0 400 80
rect 600 20 780 40
rect 600 -140 620 20
rect 760 -140 780 20
rect 600 -160 780 -140
rect 840 20 1020 40
rect 840 -140 860 20
rect 1000 -140 1020 20
rect 840 -160 1020 -140
rect 600 -240 1020 -220
rect 600 -400 660 -240
rect 960 -400 1020 -240
rect -200 -420 540 -400
rect 600 -420 1020 -400
rect -200 -580 220 -420
rect 520 -460 540 -420
rect 520 -520 860 -460
rect 520 -580 540 -520
rect -200 -600 540 -580
rect 840 -580 1020 -560
rect 600 -820 780 -600
rect 840 -740 860 -580
rect 1000 -740 1020 -580
rect 840 -760 1020 -740
rect 600 -840 1000 -820
rect 600 -900 660 -840
rect 960 -900 1000 -840
rect 600 -1000 1000 -900
rect -200 -1200 1000 -1000
<< via1 >>
rect 620 1260 760 1400
rect 620 640 760 800
rect 220 420 520 580
rect 1020 220 1180 380
rect 620 -140 760 20
rect 860 -140 1000 20
rect 220 -580 520 -420
rect 860 -740 1000 -580
<< metal2 >>
rect 600 1400 780 1420
rect 600 1260 620 1400
rect 760 1260 780 1400
rect 600 800 780 1260
rect 600 640 620 800
rect 760 640 780 800
rect 200 580 540 600
rect 200 420 220 580
rect 520 420 540 580
rect 200 400 540 420
rect 300 -400 540 400
rect 600 400 780 640
rect 600 380 1200 400
rect 600 220 1020 380
rect 1180 220 1200 380
rect 600 200 1200 220
rect 600 20 780 200
rect 600 -140 620 20
rect 760 -140 780 20
rect 600 -160 780 -140
rect 840 20 1020 40
rect 840 -140 860 20
rect 1000 -140 1020 20
rect 200 -420 540 -400
rect 200 -580 220 -420
rect 520 -580 540 -420
rect 200 -600 540 -580
rect 840 -580 1020 -140
rect 840 -740 860 -580
rect 1000 -740 1020 -580
rect 840 -760 1020 -740
use sky130_fd_pr__nfet_01v8_64Z3AY  sky130_fd_pr__nfet_01v8_64Z3AY_0 ~/tt_analog_z2a_2/mag
timestamp 1770560933
transform 1 0 811 0 1 -21
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_LGS3BL  sky130_fd_pr__pfet_01v8_LGS3BL_0 ~/tt_analog_z2a_2/mag
timestamp 1770560933
transform 1 0 811 0 1 1284
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM0
timestamp 1770560933
transform 1 0 811 0 1 -621
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_LGS3BL  XM12
timestamp 1770560933
transform 1 0 811 0 1 684
box -211 -284 211 284
<< labels >>
flabel metal1 400 -1200 600 -1000 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 400 1600 600 1800 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 200 -600 400 -400 0 FreeSans 256 0 0 0 NAND_IN_0
port 4 nsew
flabel metal1 1000 200 1200 400 0 FreeSans 256 0 0 0 NAND_OUT
port 0 nsew
flabel metal1 200 0 400 200 0 FreeSans 256 0 0 0 NAND_IN_1
port 2 nsew
<< end >>
