magic
tech sky130A
magscale 1 2
timestamp 1769857700
<< nwell >>
rect 1000 1926 2400 4200
rect 1000 1800 2362 1926
<< pwell >>
rect 1520 -1060 1900 -580
rect 1400 -1240 2000 -1060
<< viali >>
rect 1220 4100 1600 4160
rect 1820 4100 2200 4160
rect 1540 3200 1620 3880
rect 1800 3200 1880 3880
rect 1540 -800 1600 -600
rect 1820 -800 1880 -600
rect 1520 -1220 1860 -1160
rect 1920 -1920 1980 -1420
rect 1440 -2280 1940 -2240
<< metal1 >>
rect 1200 4160 2240 4600
rect 1200 4100 1220 4160
rect 1600 4100 1820 4160
rect 2200 4100 2240 4160
rect 1200 4080 2240 4100
rect 1220 3980 2060 4040
rect 1240 3340 1380 3980
rect 1520 3920 1980 3940
rect 1440 3880 1980 3920
rect 1440 3200 1540 3880
rect 1620 3200 1800 3880
rect 1880 3200 1980 3880
rect 1440 3180 1900 3200
rect 1240 840 1380 2040
rect 2040 1800 2180 2060
rect 2000 1600 2600 1800
rect 1460 1000 1980 1060
rect 1460 -200 1500 1000
rect 1920 -200 1980 1000
rect 2040 980 2180 1600
rect 1460 -240 1980 -200
rect 1520 -600 1900 -580
rect 800 -620 1200 -600
rect 800 -680 1440 -620
rect 800 -800 1200 -680
rect 1520 -800 1540 -600
rect 1600 -800 1820 -600
rect 1880 -800 1900 -600
rect 2200 -620 2600 -600
rect 1980 -680 2600 -620
rect 2200 -800 2600 -680
rect 1520 -1060 1900 -800
rect 1400 -1160 2000 -1060
rect 1400 -1220 1520 -1160
rect 1860 -1220 2000 -1160
rect 1400 -1240 2000 -1220
rect 1480 -1340 1580 -1320
rect 1200 -2120 1400 -1600
rect 1480 -2060 1500 -1340
rect 1560 -2060 1580 -1340
rect 1820 -1420 2000 -1380
rect 1820 -1920 1920 -1420
rect 1980 -1920 2000 -1420
rect 1820 -1960 2000 -1920
rect 1480 -2080 1580 -2060
rect 1200 -2180 1840 -2120
rect 1400 -2240 2000 -2220
rect 1400 -2280 1440 -2240
rect 1940 -2280 2000 -2240
rect 1400 -2600 2000 -2280
<< via1 >>
rect 1500 -200 1920 1000
rect 1500 -2060 1560 -1340
<< metal2 >>
rect 1460 1000 1980 1060
rect 1460 -200 1500 1000
rect 1920 -200 1980 1000
rect 1460 -240 1980 -200
rect 1480 -1340 1980 -240
rect 1480 -2060 1500 -1340
rect 1560 -2060 1980 -1340
rect 1480 -2080 1980 -2060
use sky130_fd_pr__nfet_01v8_A5WNKR  sky130_fd_pr__nfet_01v8_A5WNKR_0
timestamp 1768764364
transform 1 0 2011 0 1 379
box -211 -1179 211 1179
use sky130_fd_pr__pfet_01v8_MGA8MK  sky130_fd_pr__pfet_01v8_MGA8MK_0
timestamp 1769857700
transform 1 0 1411 0 1 2984
box -211 -1184 211 1184
use sky130_fd_pr__pfet_01v8_MGA8MK  XM1
timestamp 1769857700
transform 1 0 2011 0 1 2984
box -211 -1184 211 1184
use sky130_fd_pr__nfet_01v8_5ZS3RT  XM2
timestamp 1768762419
transform 1 0 1696 0 1 -1721
box -296 -579 296 579
use sky130_fd_pr__nfet_01v8_A5WNKR  XM5
timestamp 1768764364
transform 1 0 1411 0 1 379
box -211 -1179 211 1179
<< labels >>
flabel metal1 1400 -2600 1600 -2400 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 1200 -1800 1400 -1600 0 FreeSans 256 0 0 0 NBIAS
port 5 nsew
flabel metal1 1200 4400 1400 4600 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 800 -800 1000 -600 0 FreeSans 256 0 0 0 AMP_P
port 3 nsew
flabel metal1 2400 -800 2600 -600 0 FreeSans 256 0 0 0 AMP_N
port 4 nsew
rlabel metal1 2400 1600 2600 1800 1 amp_out
port 6 n default output
<< end >>
