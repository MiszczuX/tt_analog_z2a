** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/OSC5.sch
.subckt OSC5 VDD VSS OUT_OSC5
*.PININFO VDD:B VSS:B OUT_OSC5:B
x7 VDD VSS net1 OUT_OSC5 inv_x4
x9 VDD VSS net2 net1 inv_x4
x10 VDD VSS net3 net2 inv_x4
x11 VDD VSS net4 net3 inv_x4
x12 VDD VSS OUT_OSC5 net4 inv_x4
.ends

* expanding   symbol:  inv_x4.sym # of pins=4
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/inv_x4.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/inv_x4.sch
.subckt inv_x4 VDD VSS INV_OUT INV_IN
*.PININFO INV_IN:I INV_OUT:O VDD:B VSS:B
XM3 INV_OUT INV_IN VDD VDD sky130_fd_pr__pfet_01v8 L=10 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 INV_OUT INV_IN VSS VSS sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
