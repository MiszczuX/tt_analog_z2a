magic
tech sky130A
magscale 1 2
timestamp 1770560933
<< viali >>
rect 2400 -1480 2480 -1160
rect 4720 -1480 4800 -1160
rect 5200 -1480 5280 -1160
rect 7520 -1480 7600 -1160
rect 8000 -1480 8080 -1160
rect 10320 -1480 10400 -1160
rect 10800 -1480 10880 -1160
rect 13120 -1480 13200 -1160
<< metal1 >>
rect 800 800 1000 1000
rect 0 300 600 400
rect 0 -100 100 300
rect 500 200 600 300
rect 14600 300 15200 400
rect 500 0 800 200
rect 500 -100 600 0
rect 0 -200 600 -100
rect 14600 -100 14700 300
rect 15100 -100 15200 300
rect 14600 -200 15200 -100
rect 800 -400 1000 -200
rect 2300 -1160 2500 -700
rect 2300 -1480 2400 -1160
rect 2480 -1300 2500 -1160
rect 3400 -1020 3800 -1000
rect 3400 -1180 3420 -1020
rect 3780 -1180 3800 -1020
rect 3400 -1200 3800 -1180
rect 4700 -1160 5300 -800
rect 4700 -1300 4720 -1160
rect 2480 -1480 2600 -1300
rect 2300 -1600 2600 -1480
rect 4600 -1480 4720 -1300
rect 4800 -1480 5200 -1160
rect 5280 -1300 5300 -1160
rect 6200 -1020 6600 -1000
rect 6200 -1180 6220 -1020
rect 6580 -1180 6600 -1020
rect 6200 -1200 6600 -1180
rect 7500 -1160 8100 -700
rect 10700 -800 10900 -700
rect 7500 -1300 7520 -1160
rect 5280 -1480 5400 -1300
rect 4600 -1600 5400 -1480
rect 7400 -1480 7520 -1300
rect 7600 -1480 8000 -1160
rect 8080 -1300 8100 -1160
rect 9000 -1020 9400 -1000
rect 9000 -1180 9020 -1020
rect 9380 -1180 9400 -1020
rect 9000 -1200 9400 -1180
rect 10300 -1160 10900 -800
rect 10300 -1300 10320 -1160
rect 8080 -1480 8200 -1300
rect 7400 -1600 8200 -1480
rect 10200 -1480 10320 -1300
rect 10400 -1480 10800 -1160
rect 10880 -1300 10900 -1160
rect 11800 -1020 12200 -1000
rect 11800 -1180 11820 -1020
rect 12180 -1180 12200 -1020
rect 11800 -1200 12200 -1180
rect 13100 -1160 13300 -700
rect 13100 -1300 13120 -1160
rect 10880 -1480 11000 -1300
rect 10200 -1600 11000 -1480
rect 13000 -1480 13120 -1300
rect 13200 -1480 13300 -1160
rect 13000 -1600 13300 -1480
<< via1 >>
rect 100 -100 500 300
rect 3420 20 3780 180
rect 6220 20 6580 180
rect 9020 20 9380 180
rect 11820 20 12180 180
rect 14700 -100 15100 300
rect 3420 -1180 3780 -1020
rect 6220 -1180 6580 -1020
rect 9020 -1180 9380 -1020
rect 11820 -1180 12180 -1020
<< metal2 >>
rect 0 600 15200 1000
rect 0 300 600 600
rect 0 -100 100 300
rect 500 -100 600 300
rect 14600 300 15200 600
rect 0 -200 600 -100
rect 3400 180 3800 200
rect 3400 20 3420 180
rect 3780 20 3800 180
rect 3400 -1020 3800 20
rect 3400 -1180 3420 -1020
rect 3780 -1180 3800 -1020
rect 3400 -1200 3800 -1180
rect 6200 180 6600 200
rect 6200 20 6220 180
rect 6580 20 6600 180
rect 6200 -1020 6600 20
rect 6200 -1180 6220 -1020
rect 6580 -1180 6600 -1020
rect 6200 -1200 6600 -1180
rect 9000 180 9400 200
rect 9000 20 9020 180
rect 9380 20 9400 180
rect 9000 -1020 9400 20
rect 9000 -1180 9020 -1020
rect 9380 -1180 9400 -1020
rect 9000 -1200 9400 -1180
rect 11800 180 12200 200
rect 11800 20 11820 180
rect 12180 20 12200 180
rect 11800 -1020 12200 20
rect 14600 -100 14700 300
rect 15100 -100 15200 300
rect 14600 -200 15200 -100
rect 11800 -1180 11820 -1020
rect 12180 -1180 12200 -1020
rect 11800 -1200 12200 -1180
use sky130_fd_pr__nfet_01v8_QXQT3M  sky130_fd_pr__nfet_01v8_QXQT3M_0 ~/tt_analog_z2a_2/mag
timestamp 1770560933
transform 1 0 11997 0 1 -1320
box -1196 -279 1196 279
use inv_x4  x22 ~/tt_analog_z2a_2/mag
timestamp 1770560933
transform 1 0 0 0 1 400
box 800 -1200 3600 800
use inv_x4  x23
timestamp 1770560933
transform 1 0 2800 0 1 400
box 800 -1200 3600 800
use inv_x4  x24
timestamp 1770560933
transform 1 0 5600 0 1 400
box 800 -1200 3600 800
use inv_x4  x25
timestamp 1770560933
transform 1 0 8400 0 1 400
box 800 -1200 3600 800
use inv_x4  x26
timestamp 1770560933
transform 1 0 11200 0 1 400
box 800 -1200 3600 800
use sky130_fd_pr__nfet_01v8_QXQT3M  XM1
timestamp 1770560933
transform 1 0 6397 0 1 -1320
box -1196 -279 1196 279
use sky130_fd_pr__nfet_01v8_QXQT3M  XM2
timestamp 1770560933
transform 1 0 9197 0 1 -1320
box -1196 -279 1196 279
use sky130_fd_pr__nfet_01v8_QXQT3M  XM5
timestamp 1770560933
transform 1 0 3597 0 1 -1320
box -1196 -279 1196 279
<< labels >>
flabel metal1 800 800 1000 1000 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 800 -400 1000 -200 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel via1 14800 0 15000 200 0 FreeSans 256 0 0 0 OUT_OSC5cap
port 2 nsew
<< end >>
