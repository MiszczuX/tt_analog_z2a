** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/OSC3.sch
.subckt OSC3 VDD VSS OUT_OSC3
*.PININFO VDD:B VSS:B OUT_OSC3:B
x19 VDD VSS net1 OUT_OSC3 inv_x4
x20 VDD VSS net2 net1 inv_x4
x21 VDD VSS OUT_OSC3 net2 inv_x4
.ends

* expanding   symbol:  inv_x4.sym # of pins=4
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/inv_x4.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/inv_x4.sch
.subckt inv_x4 VDD VSS INV_OUT INV_IN
*.PININFO INV_IN:I INV_OUT:O VDD:B VSS:B
XM3 INV_OUT INV_IN VDD VDD sky130_fd_pr__pfet_01v8 L=10 W=2 nf=1 m=1
XM5 INV_OUT INV_IN VSS VSS sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
.ends

.end
