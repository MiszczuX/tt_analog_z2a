magic
tech sky130A
timestamp 1768677564
<< metal1 >>
rect -2238 1743 -700 1800
rect -2249 1700 -700 1743
rect -2249 -213 -2086 1700
rect -1400 1300 -800 1400
rect 3100 900 4000 1000
rect -1450 650 -1350 700
rect -1450 640 -1000 650
rect -1450 610 -1090 640
rect -1010 610 -1000 640
rect -1450 600 -1000 610
rect -1600 550 -1500 600
rect -1600 540 -900 550
rect -1600 510 -990 540
rect -910 510 -900 540
rect -1600 500 -900 510
rect -1750 450 -1650 500
rect -1750 440 -800 450
rect -1750 410 -890 440
rect -810 410 -800 440
rect -1750 400 -800 410
rect -1900 350 -1800 400
rect -1900 340 -700 350
rect -1900 310 -790 340
rect -710 310 -700 340
rect -1900 300 -700 310
rect -1800 240 -600 250
rect -1800 210 -690 240
rect -610 210 -600 240
rect -1800 200 -600 210
rect -1800 150 -1700 200
rect -1650 140 -500 150
rect -1650 110 -590 140
rect -510 110 -500 140
rect -1650 100 -500 110
rect 3900 100 4000 900
rect -1650 50 -1550 100
rect -1500 40 -430 50
rect -1500 10 -490 40
rect -440 10 -430 40
rect -1500 0 -430 10
rect 3500 0 4000 100
rect -1500 -50 -1400 0
rect -2249 -346 -1506 -213
rect -2249 -393 -1764 -346
rect -1611 -393 -1506 -346
rect -2249 -467 -1506 -393
rect -1200 -1362 -1150 -250
rect -1100 -1348 -1050 -250
rect -1000 -1264 -950 -250
rect -900 -1187 -850 -250
rect -800 -1152 -750 -250
rect -1209 -2535 -1139 -1362
rect -1111 -2521 -1041 -1348
rect -1006 -2437 -936 -1264
rect -902 -2360 -832 -1187
rect -811 -2325 -741 -1152
rect -1200 -2660 -1150 -2535
rect -1200 -2740 -1190 -2660
rect -1160 -2740 -1150 -2660
rect -1200 -3105 -1150 -2740
rect -1100 -3105 -1050 -2521
rect -1000 -3105 -950 -2437
rect -900 -3105 -850 -2360
rect -800 -3105 -750 -2325
rect -700 -3105 -650 -250
rect -600 -3105 -550 -250
rect -500 -3105 -450 -250
rect -400 -3105 -350 -100
rect -300 -2360 -250 -150
rect -300 -2440 -290 -2360
rect -260 -2440 -250 -2360
rect -300 -3105 -250 -2440
rect -200 -2060 -150 -150
rect -200 -2140 -190 -2060
rect -160 -2140 -150 -2060
rect -200 -3105 -150 -2140
rect -100 -1760 -50 -150
rect -100 -1840 -90 -1760
rect -60 -1840 -50 -1760
rect -100 -3105 -50 -1840
rect 0 -1460 50 -150
rect 0 -1540 10 -1460
rect 40 -1540 50 -1460
rect 0 -3105 50 -1540
rect 100 -1160 150 -150
rect 100 -1240 110 -1160
rect 140 -1240 150 -1160
rect 100 -3105 150 -1240
rect 200 -860 250 -150
rect 200 -940 210 -860
rect 240 -940 250 -860
rect 200 -3105 250 -940
rect 300 -560 350 -150
rect 500 -400 600 -300
rect 1600 -400 1800 -300
rect 300 -640 310 -560
rect 340 -640 350 -560
rect 300 -3105 350 -640
rect 1900 -1700 2000 -1600
rect 400 -2450 500 -2400
rect 1451 -3193 1600 -3079
rect 1800 -3079 1900 -2000
rect 1800 -3193 1954 -3079
rect 1451 -3289 1954 -3193
<< via1 >>
rect -690 1310 -610 1390
rect -1090 610 -1010 640
rect -990 510 -910 540
rect -890 410 -810 440
rect -790 310 -710 340
rect -690 210 -610 240
rect -590 110 -510 140
rect 3500 100 3900 900
rect -490 10 -440 40
rect -1764 -393 -1611 -346
rect -1190 -2740 -1160 -2660
rect -290 -2440 -260 -2360
rect -190 -2140 -160 -2060
rect -90 -1840 -60 -1760
rect 10 -1540 40 -1460
rect 110 -1240 140 -1160
rect 210 -940 240 -860
rect 310 -640 340 -560
rect 1600 -3193 1800 -2100
<< metal2 >>
rect 3400 900 4000 1000
rect 3900 100 4000 900
rect -1824 -313 -1544 -293
rect -1251 -313 600 -300
rect -1824 -346 600 -313
rect -1824 -393 -1764 -346
rect -1611 -393 600 -346
rect -1824 -400 600 -393
rect -1824 -420 -1192 -400
rect -1824 -453 -1544 -420
rect -1251 -560 700 -550
rect -1251 -640 310 -560
rect 340 -640 700 -560
rect -1251 -650 700 -640
rect -1251 -860 700 -850
rect -1251 -940 210 -860
rect 240 -940 700 -860
rect -1251 -950 700 -940
rect -1244 -1160 700 -1150
rect -1244 -1240 110 -1160
rect 140 -1240 700 -1160
rect -1244 -1250 700 -1240
rect 0 -1460 700 -1450
rect 0 -1540 10 -1460
rect 40 -1540 700 -1460
rect 0 -1550 700 -1540
rect -100 -1760 700 -1750
rect -100 -1840 -90 -1760
rect -60 -1840 700 -1760
rect -100 -1850 700 -1840
rect 3500 -2000 4000 100
rect -200 -2060 700 -2050
rect -200 -2140 -190 -2060
rect -160 -2140 700 -2060
rect -200 -2150 700 -2140
rect 1500 -2100 4000 -2000
rect -300 -2360 700 -2350
rect -300 -2440 -290 -2360
rect -260 -2440 700 -2360
rect -300 -2450 700 -2440
rect -1244 -2660 700 -2650
rect -1244 -2740 -1190 -2660
rect -1160 -2740 700 -2660
rect -1244 -2750 700 -2740
rect -1244 -3100 500 -2900
rect 1500 -3079 1600 -2100
rect 1451 -3193 1600 -3079
rect 1800 -3000 4000 -2100
rect 1800 -3079 1900 -3000
rect 1800 -3193 1954 -3079
rect 1451 -3289 1954 -3193
use AND  x1
timestamp 1768672672
transform 1 0 450 0 1 -750
box 50 -2250 1550 450
use LOGIC_INV  x9
timestamp 1768674023
transform 1 0 -1000 0 1 4600
box -200 -4850 4300 -2700
<< labels >>
flabel metal1 500 -400 600 -300 0 FreeSans 128 0 0 0 VDD
port 17 nsew
flabel metal1 1900 -1700 2000 -1600 0 FreeSans 128 0 0 0 LOGICOUT_0_2
port 16 nsew
flabel metal1 -1350 1300 -1250 1400 0 FreeSans 128 0 0 0 LOGICIN_0_2
port 12 nsew
flabel metal1 -1450 600 -1350 700 0 FreeSans 128 0 0 0 LOGICIN_0_4
port 11 nsew
flabel metal1 -1600 500 -1500 600 0 FreeSans 128 0 0 0 LOGICIN_0_6
port 10 nsew
flabel metal1 -1750 400 -1650 500 0 FreeSans 128 0 0 0 LOGICIN_0_8
port 8 nsew
flabel metal1 -1900 300 -1800 400 0 FreeSans 128 0 0 0 LOGICIN_1_0
port 7 nsew
flabel metal1 -1800 150 -1700 250 0 FreeSans 128 0 0 0 LOGICIN_1_2
port 6 nsew
flabel metal1 -1650 50 -1550 150 0 FreeSans 128 0 0 0 LOGICIN_1_4
port 5 nsew
flabel metal1 -1500 -50 -1400 50 0 FreeSans 128 0 0 0 LOGICIN_1_6
port 4 nsew
<< end >>
