** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/yen_top.sch
.subckt yen_top VDD VSS VCMUXIN VCMUXOUT
*.PININFO VDD:B VSS:B VCMUXIN:B VCMUXOUT:B
x2 vbg_1_6 vbg_1_4 vbg_1_2 vbg_1_0 vbg_0_8 vbg_0_6 vbg_0_4 vbg_0_2 VDD VSS BG
x1 in_1_6 VCMUXOUT in_1_4 in_1_2 in_1_0 in_0_8 in_0_6 in_0_4 in_0_2 vbg_1_6 VDD vbg_1_4 VSS vbg_1_2 vbg_1_0 vbg_0_8 vbg_0_6
+ vbg_0_4 vbg_0_2 VCMUXIN VCMUX
x5 in_0_8 VDD in_0_6 in_0_4 VDD VSS T_FLIP_FLOP
x7 VDD VSS in_1_2 in_1_0 inv_x1
x9 bg16 bg14 bg12 bg10 bg08 bg06 bg04 in_1_6 VDD VSS BG
x3 VDD VSS in_0_2 OSC3
x4 VDD VSS in_0_6 OSC5
x6 VDD VSS in_1_0 OSC7
x8 VDD VSS in_1_4 OSC5cap
.ends

* expanding   symbol:  BG.sym # of pins=10
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/BG.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/BG.sch
.subckt BG vbg_1_6 vbg_1_4 vbg_1_2 vbg_1_0 vbg_0_8 vbg_0_6 vbg_0_4 vbg_0_2 VDD VSS
*.PININFO vbg_1_6:O vbg_1_4:O vbg_1_2:O vbg_1_0:O vbg_0_8:O vbg_0_6:O vbg_0_4:O vbg_0_2:O VDD:B VSS:B
XR1 vbg_1_4 vbg_1_6 VSS sky130_fd_pr__res_high_po_0p35 L=1.5 mult=1 m=1
XR0 vbg_1_6 VDD VSS sky130_fd_pr__res_high_po_0p35 L=1.5 mult=1 m=1
XR3 vbg_1_0 vbg_1_2 VSS sky130_fd_pr__res_high_po_0p35 L=1.5 mult=1 m=1
XR2 vbg_1_2 vbg_1_4 VSS sky130_fd_pr__res_high_po_0p35 L=1.5 mult=1 m=1
XR5 vbg_0_6 vbg_0_8 VSS sky130_fd_pr__res_high_po_0p35 L=1.5 mult=1 m=1
XR4 vbg_0_8 vbg_1_0 VSS sky130_fd_pr__res_high_po_0p35 L=1.5 mult=1 m=1
XR6 vbg_0_4 vbg_0_6 VSS sky130_fd_pr__res_high_po_0p35 L=1.5 mult=1 m=1
XR7 vbg_0_2 vbg_0_4 VSS sky130_fd_pr__res_high_po_0p35 L=1.5 mult=1 m=1
XR8 VSS vbg_0_2 VSS sky130_fd_pr__res_high_po_0p35 L=1.5 mult=1 m=1
.ends


* expanding   symbol:  VCMUX.sym # of pins=20
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/VCMUX.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/VCMUX.sch
.subckt VCMUX VCMUX_IN_1_6 VCMUX_OUT VCMUX_IN_1_4 VCMUX_IN_1_2 VCMUX_IN_1_0 VCMUX_IN_0_8 VCMUX_IN_0_6 VCMUX_IN_0_4 VCMUX_IN_0_2
+ vbg_1_6 VDD vbg_1_4 VSS vbg_1_2 vbg_1_0 vbg_0_8 vbg_0_6 vbg_0_4 vbg_0_2 VCMUX_IN
*.PININFO VDD:B VSS:B vbg_1_6:I vbg_1_4:I vbg_1_2:I vbg_1_0:I vbg_0_8:I vbg_0_6:I vbg_0_4:I vbg_0_2:I VCMUX_IN:I VCMUX_IN_0_2:I
*+ VCMUX_IN_0_4:I VCMUX_IN_0_6:I VCMUX_IN_0_8:I VCMUX_IN_1_0:I VCMUX_IN_1_2:I VCMUX_OUT:O VCMUX_IN_1_4:I VCMUX_IN_1_6:I
x0 VDD VSS vbg_0_6 VCMUX_IN DISC_OUT_0_2 vbg_0_2 pdiscr
x1 VDD VSS vbg_0_6 VCMUX_IN DISC_OUT_0_4 vbg_0_4 pdiscr
x2 VDD VSS vbg_0_6 VCMUX_IN DISC_OUT_0_6 vbg_0_6 pdiscr
x3 VDD VSS vbg_0_6 VCMUX_IN DISC_OUT_0_8 vbg_0_8 pdiscr
x4 VDD VSS vbg_1_0 VCMUX_IN DISC_OUT_1_0 vbg_1_0 ndiscr
x5 VDD VSS vbg_1_0 VCMUX_IN DISC_OUT_1_2 vbg_1_2 ndiscr
x6 VDD VSS vbg_1_0 VCMUX_IN DISC_OUT_1_4 vbg_1_4 ndiscr
x7 VDD VSS vbg_1_0 VCMUX_IN DISC_OUT_1_6 vbg_1_6 ndiscr
x8 LOGIC_OUT_1_6 LOGIC_OUT_1_4 LOGIC_OUT_1_2 LOGIC_OUT_1_0 DISC_OUT_1_6 DISC_OUT_1_4 DISC_OUT_1_2 DISC_OUT_1_0 DISC_OUT_0_8
+ DISC_OUT_0_6 DISC_OUT_0_4 DISC_OUT_0_2 LOGIC_OUT_0_8 LOGIC_OUT_0_6 LOGIC_OUT_0_4 LOGIC_OUT_0_2 VDD VSS LOGIC
x9 VDD VCMUX_IN_0_2 VSS LOGIC_OUT_0_2 VCMUX_OUT PASSGATE
x10 VDD VCMUX_IN_0_4 VSS LOGIC_OUT_0_4 VCMUX_OUT PASSGATE
x11 VDD VCMUX_IN_0_6 VSS LOGIC_OUT_0_6 VCMUX_OUT PASSGATE
x12 VDD VCMUX_IN_0_8 VSS LOGIC_OUT_0_8 VCMUX_OUT PASSGATE
x13 VDD VCMUX_IN_1_0 VSS LOGIC_OUT_1_0 VCMUX_OUT PASSGATE
x14 VDD VCMUX_IN_1_2 VSS LOGIC_OUT_1_2 VCMUX_OUT PASSGATE
x15 VDD VCMUX_IN_1_4 VSS LOGIC_OUT_1_4 VCMUX_OUT PASSGATE
x16 VDD VCMUX_IN_1_6 VSS LOGIC_OUT_1_6 VCMUX_OUT PASSGATE
.ends


* expanding   symbol:  T_FLIP_FLOP.sym # of pins=6
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/T_FLIP_FLOP.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/T_FLIP_FLOP.sch
.subckt T_FLIP_FLOP Q T_IN CLK ZQ VDD VSS
*.PININFO VDD:B VSS:B CLK:I ZQ:O Q:O T_IN:I
x2 ZQ VDD out1 VSS Q NAND2
x4 Q VDD out2 VSS ZQ NAND2
x1 out1 VDD CLK VSS net1 NAND2
x3 out2 VDD T_IN VSS CLK NAND2
x24 VDD VSS net1 T_IN inv_x4
.ends


* expanding   symbol:  inv_x1.sym # of pins=4
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/inv_x1.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/inv_x1.sch
.subckt inv_x1 VDD VSS INV_OUT INV_IN
*.PININFO INV_IN:I INV_OUT:O VDD:B VSS:B
XM3 INV_OUT INV_IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 INV_OUT INV_IN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  OSC3.sym # of pins=3
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/OSC3.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/OSC3.sch
.subckt OSC3 VDD VSS OUT_OSC3
*.PININFO VDD:B VSS:B OUT_OSC3:B
x19 VDD VSS net1 OUT_OSC3 inv_x4
x20 VDD VSS net2 net1 inv_x4
x21 VDD VSS OUT_OSC3 net2 inv_x4
.ends


* expanding   symbol:  OSC5.sym # of pins=3
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/OSC5.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/OSC5.sch
.subckt OSC5 VDD VSS OUT_OSC5
*.PININFO VDD:B VSS:B OUT_OSC5:B
x7 VDD VSS net1 OUT_OSC5 inv_x4
x9 VDD VSS net2 net1 inv_x4
x10 VDD VSS net3 net2 inv_x4
x11 VDD VSS net4 net3 inv_x4
x12 VDD VSS OUT_OSC5 net4 inv_x4
.ends


* expanding   symbol:  OSC7.sym # of pins=3
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/OSC7.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/OSC7.sch
.subckt OSC7 VDD VSS OUT_OSC7
*.PININFO VDD:B VSS:B OUT_OSC7:B
x8 VDD VSS net1 OUT_OSC7 inv_x4
x5 VDD VSS net2 net1 inv_x4
x6 VDD VSS net3 net2 inv_x4
x13 VDD VSS net4 net3 inv_x4
x14 VDD VSS net5 net4 inv_x4
x15 VDD VSS net6 net5 inv_x4
x16 VDD VSS OUT_OSC7 net6 inv_x4
.ends


* expanding   symbol:  OSC5cap.sym # of pins=3
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/OSC5cap.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/OSC5cap.sch
.subckt OSC5cap VDD VSS OUT_OSC5cap
*.PININFO VDD:B VSS:B OUT_OSC5cap:B
x22 VDD VSS net1 OUT_OSC5cap inv_x4
x23 VDD VSS net2 net1 inv_x4
x24 VDD VSS net3 net2 inv_x4
x25 VDD VSS net4 net3 inv_x4
x26 VDD VSS OUT_OSC5cap net4 inv_x4
XM5 VSS net1 VSS VSS sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
XM1 VSS net2 VSS VSS sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
XM2 VSS net3 VSS VSS sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
XM3 VSS net4 VSS VSS sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
.ends


* expanding   symbol:  pdiscr.sym # of pins=6
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/pdiscr.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/pdiscr.sch
.subckt pdiscr VDD VSS DISCR_BIAS DISCR_IN DISCR_OUT DISCR_VREF
*.PININFO VDD:B VSS:B DISCR_IN:I DISCR_VREF:I DISCR_OUT:O DISCR_BIAS:B
x6 VDD VSS net2 net1 inv_x1
x7 VDD VSS DISCR_OUT net2 inv_x1
x5 VDD VSS net1 DISCR_IN DISCR_VREF DISCR_BIAS amp_p
.ends


* expanding   symbol:  ndiscr.sym # of pins=6
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/ndiscr.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/ndiscr.sch
.subckt ndiscr VDD VSS DISCR_BIAS DISCR_IN DISCR_OUT DISCR_VREF
*.PININFO VDD:B VSS:B DISCR_IN:I DISCR_VREF:I DISCR_OUT:O DISCR_BIAS:B
x6 VDD VSS net2 net1 inv_x1
x7 VDD VSS DISCR_OUT net2 inv_x1
x17 VDD VSS net1 DISCR_IN DISCR_VREF DISCR_BIAS amp
.ends


* expanding   symbol:  LOGIC.sym # of pins=18
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/LOGIC.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/LOGIC.sch
.subckt LOGIC LOGICOUT_1_6 LOGICOUT_1_4 LOGICOUT_1_2 LOGICOUT_1_0 LOGICIN_1_6 LOGICIN_1_4 LOGICIN_1_2 LOGICIN_1_0 LOGICIN_0_8
+ LOGICIN_0_6 LOGICIN_0_4 LOGICIN_0_2 LOGICOUT_0_8 LOGICOUT_0_6 LOGICOUT_0_4 LOGICOUT_0_2 VDD VSS
*.PININFO LOGICOUT_0_2:O LOGICOUT_0_4:O LOGICOUT_0_6:O LOGICOUT_0_8:O LOGICOUT_1_0:O LOGICOUT_1_2:O LOGICOUT_1_4:O LOGICOUT_1_6:O
*+ LOGICIN_1_0:I LOGICIN_1_2:I LOGICIN_1_4:I LOGICIN_1_6:I LOGICIN_0_2:I LOGICIN_0_4:I LOGICIN_0_6:I LOGICIN_0_8:I VDD:B VSS:B
x1 VDD VSS Z_LOGICIN_1_6 Z_LOGICIN_1_4 Z_LOGICIN_1_2 Z_LOGICIN_1_0 LOGICOUT_0_2 Z_LOGICIN_0_8 Z_LOGICIN_0_6 Z_LOGICIN_0_4
+ LOGICIN_0_2 AND
x2 VDD VSS Z_LOGICIN_1_6 Z_LOGICIN_1_4 Z_LOGICIN_1_2 Z_LOGICIN_1_0 LOGICOUT_0_4 Z_LOGICIN_0_8 Z_LOGICIN_0_6 LOGICIN_0_4
+ LOGICIN_0_2 AND
x3 VDD VSS Z_LOGICIN_1_6 Z_LOGICIN_1_4 Z_LOGICIN_1_2 Z_LOGICIN_1_0 LOGICOUT_0_6 Z_LOGICIN_0_8 LOGICIN_0_6 LOGICIN_0_4 LOGICIN_0_2
+ AND
x4 VDD VSS Z_LOGICIN_1_6 Z_LOGICIN_1_4 Z_LOGICIN_1_2 Z_LOGICIN_1_0 LOGICOUT_0_8 LOGICIN_0_8 LOGICIN_0_6 LOGICIN_0_4 LOGICIN_0_2
+ AND
x5 VDD VSS Z_LOGICIN_1_6 Z_LOGICIN_1_4 Z_LOGICIN_1_2 LOGICIN_1_0 LOGICOUT_1_0 LOGICIN_0_8 LOGICIN_0_6 LOGICIN_0_4 LOGICIN_0_2 AND
x6 VDD VSS Z_LOGICIN_1_6 Z_LOGICIN_1_4 LOGICIN_1_2 LOGICIN_1_0 LOGICOUT_1_2 LOGICIN_0_8 LOGICIN_0_6 LOGICIN_0_4 LOGICIN_0_2 AND
x7 VDD VSS Z_LOGICIN_1_6 LOGICIN_1_4 LOGICIN_1_2 LOGICIN_1_0 LOGICOUT_1_4 LOGICIN_0_8 LOGICIN_0_6 LOGICIN_0_4 LOGICIN_0_2 AND
x8 VDD VSS LOGICIN_1_6 LOGICIN_1_4 LOGICIN_1_2 LOGICIN_1_0 LOGICOUT_1_6 LOGICIN_0_8 LOGICIN_0_6 LOGICIN_0_4 LOGICIN_0_2 AND
x9 LOGICIN_1_6 Z_LOGICIN_1_6 Z_LOGICIN_1_4 LOGICIN_1_4 LOGICIN_1_2 Z_LOGICIN_1_2 LOGICIN_1_0 Z_LOGICIN_1_0 Z_LOGICIN_0_8
+ LOGICIN_0_8 Z_LOGICIN_0_6 LOGICIN_0_6 LOGICIN_0_4 Z_LOGICIN_0_4 LOGICIN_0_2 Z_LOGICIN_0_2 VDD VSS LOGIC_INV
.ends


* expanding   symbol:  PASSGATE.sym # of pins=5
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/PASSGATE.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/PASSGATE.sch
.subckt PASSGATE VDD PASS_GATE_IN VSS PASS_GATE_EN PASS_GATE_OUT
*.PININFO PASS_GATE_IN:B PASS_GATE_EN:I VDD:B VSS:B PASS_GATE_OUT:B
XM1pass PASS_GATE_ZEN PASS_GATE_EN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=10 nf=1 m=1
XM0pass PASS_GATE_ZEN PASS_GATE_EN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 m=1
XM1 PASS_GATE_IN PASS_GATE_EN PASS_GATE_OUT VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 PASS_GATE_OUT PASS_GATE_ZEN PASS_GATE_IN VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  NAND2.sym # of pins=5
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/NAND2.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/NAND2.sch
.subckt NAND2 NAND_OUT VDD NAND_IN_1 VSS NAND_IN_0
*.PININFO NAND_IN_0:I NAND_OUT:O VDD:B VSS:B NAND_IN_1:I
XM0 net1 NAND_IN_0 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM1 NAND_OUT NAND_IN_1 net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM12 NAND_OUT NAND_IN_0 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM13 NAND_OUT NAND_IN_1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  inv_x4.sym # of pins=4
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/inv_x4.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/inv_x4.sch
.subckt inv_x4 VDD VSS INV_OUT INV_IN
*.PININFO INV_IN:I INV_OUT:O VDD:B VSS:B
XM3 INV_OUT INV_IN VDD VDD sky130_fd_pr__pfet_01v8 L=10 W=2 nf=1 m=1
XM5 INV_OUT INV_IN VSS VSS sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
.ends


* expanding   symbol:  amp_p.sym # of pins=6
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/amp_p.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/amp_p.sch
.subckt amp_p VDD VSS AMP_OUT AMP_P AMP_N PBIAS
*.PININFO AMP_P:I AMP_N:I AMP_OUT:O PBIAS:I VDD:B VSS:B
XM1 VTAIL PBIAS VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=8 nf=1 m=1
XM2 AMP_OUT VFOLD VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 m=1
XM6 VFOLD VFOLD VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 m=1
XM4 AMP_OUT AMP_N VTAIL VDD sky130_fd_pr__pfet_01v8 L=0.15 W=10 nf=2 m=1
XM5 VFOLD AMP_P VTAIL VDD sky130_fd_pr__pfet_01v8 L=0.15 W=10 nf=2 m=1
.ends


* expanding   symbol:  amp.sym # of pins=6
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/amp.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/amp.sch
.subckt amp VDD VSS AMP_OUT AMP_P AMP_N NBIAS
*.PININFO AMP_P:I AMP_N:I AMP_OUT:O NBIAS:I VDD:B VSS:B
XM3 VFOLD VFOLD VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=10 nf=1 m=1
XM4 AMP_OUT AMP_N VTAIL VSS sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 m=1
XM1 AMP_OUT VFOLD VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=10 nf=1 m=1
XM5 VFOLD AMP_P VTAIL VSS sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 m=1
XM2 VTAIL NBIAS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=4 nf=1 m=1
.ends


* expanding   symbol:  AND.sym # of pins=11
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/AND.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/AND.sch
.subckt AND VDD VSS AND_IN_1_6 AND_IN_1_4 AND_IN_1_2 AND_IN_1_0 AND_OUT AND_IN_0_8 AND_IN_0_6 AND_IN_0_4 AND_IN_0_2
*.PININFO VDD:B VSS:B AND_IN_0_2:I AND_OUT:O AND_IN_0_4:I AND_IN_0_6:I AND_IN_0_8:I AND_IN_1_0:I AND_IN_1_2:I AND_IN_1_4:I
*+ AND_IN_1_6:I
x5 NANDOUT AND_IN_1_6 VDD AND_IN_1_4 VSS AND_IN_1_2 AND_IN_1_0 AND_IN_0_8 AND_IN_0_6 AND_IN_0_4 AND_IN_0_2 NAND
x28 VDD VSS AND_OUT NANDOUT inv_x1
.ends


* expanding   symbol:  LOGIC_INV.sym # of pins=18
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/LOGIC_INV.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/LOGIC_INV.sch
.subckt LOGIC_INV LOGICIN_1_6 Z_LOGICIN_1_6 Z_LOGICIN_1_4 LOGICIN_1_4 LOGICIN_1_2 Z_LOGICIN_1_2 LOGICIN_1_0 Z_LOGICIN_1_0
+ Z_LOGICIN_0_8 LOGICIN_0_8 Z_LOGICIN_0_6 LOGICIN_0_6 LOGICIN_0_4 Z_LOGICIN_0_4 LOGICIN_0_2 Z_LOGICIN_0_2 VDD VSS
*.PININFO Z_LOGICIN_0_2:O LOGICIN_0_2:I LOGICIN_0_4:I LOGICIN_0_6:I LOGICIN_0_8:I LOGICIN_1_0:I LOGICIN_1_2:I LOGICIN_1_4:I
*+ LOGICIN_1_6:I Z_LOGICIN_0_4:O Z_LOGICIN_0_6:O Z_LOGICIN_0_8:O Z_LOGICIN_1_0:O Z_LOGICIN_1_2:O Z_LOGICIN_1_4:O Z_LOGICIN_1_6:O VDD:B VSS:B
x28 VDD VSS Z_LOGICIN_0_2 LOGICIN_0_2 inv_x1
x1 VDD VSS Z_LOGICIN_0_4 LOGICIN_0_4 inv_x1
x2 VDD VSS Z_LOGICIN_0_6 LOGICIN_0_6 inv_x1
x3 VDD VSS Z_LOGICIN_0_8 LOGICIN_0_8 inv_x1
x4 VDD VSS Z_LOGICIN_1_0 LOGICIN_1_0 inv_x1
x5 VDD VSS Z_LOGICIN_1_2 LOGICIN_1_2 inv_x1
x6 VDD VSS Z_LOGICIN_1_4 LOGICIN_1_4 inv_x1
x7 VDD VSS Z_LOGICIN_1_6 LOGICIN_1_6 inv_x1
.ends


* expanding   symbol:  NAND.sym # of pins=11
** sym_path: /home/ttuser/tt_analog_z2a_2/xschem/NAND.sym
** sch_path: /home/ttuser/tt_analog_z2a_2/xschem/NAND.sch
.subckt NAND NAND_OUT NAND_IN_7 VDD NAND_IN_6 VSS NAND_IN_5 NAND_IN_4 NAND_IN_3 NAND_IN_2 NAND_IN_1 NAND_IN_0
*.PININFO NAND_IN_0:I NAND_OUT:O VDD:B VSS:B NAND_IN_1:I NAND_IN_2:I NAND_IN_3:I NAND_IN_4:I NAND_IN_5:I NAND_IN_6:I NAND_IN_7:I
XM15 NAND_OUT NAND_IN_0 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM0 net1 NAND_IN_0 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM1 net2 NAND_IN_1 net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 net3 NAND_IN_2 net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 net4 NAND_IN_3 net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net5 NAND_IN_4 net4 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 net6 NAND_IN_5 net5 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 net7 NAND_IN_6 net6 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM7 NAND_OUT NAND_IN_7 net7 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM8 NAND_OUT NAND_IN_1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM9 NAND_OUT NAND_IN_2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM10 NAND_OUT NAND_IN_3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM11 NAND_OUT NAND_IN_4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM12 NAND_OUT NAND_IN_5 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM13 NAND_OUT NAND_IN_6 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM14 NAND_OUT NAND_IN_7 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

.end
