** sch_path: /home/ttuser/tt_analog_z2a/xschem/NAND.sch
.subckt NAND NAND_OUT NAND_IN_7 VDD NAND_IN_6 VSS NAND_IN_5 NAND_IN_4 NAND_IN_3 NAND_IN_2 NAND_IN_1 NAND_IN_0
*.PININFO NAND_IN_0:I NAND_OUT:O VDD:B VSS:B NAND_IN_1:I NAND_IN_2:I NAND_IN_3:I NAND_IN_4:I NAND_IN_5:I NAND_IN_6:I NAND_IN_7:I
XM15 NAND_OUT NAND_IN_0 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM0 net1 NAND_IN_0 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM1 net2 NAND_IN_1 net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 net3 NAND_IN_2 net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 net4 NAND_IN_3 net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net5 NAND_IN_4 net4 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 net6 NAND_IN_5 net5 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 net7 NAND_IN_6 net6 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM7 NAND_OUT NAND_IN_7 net7 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM8 NAND_OUT NAND_IN_1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM9 NAND_OUT NAND_IN_2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM10 NAND_OUT NAND_IN_3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM11 NAND_OUT NAND_IN_4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM12 NAND_OUT NAND_IN_5 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM13 NAND_OUT NAND_IN_6 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM14 NAND_OUT NAND_IN_7 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends
.end
