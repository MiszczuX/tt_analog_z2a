magic
tech sky130A
magscale 1 2
timestamp 1769862601
<< nwell >>
rect 800 -4300 1300 400
rect 800 -4400 1100 -4300
<< pwell >>
rect 380 -2100 640 -2060
rect 380 -2580 640 -2540
rect 380 -2700 640 -2660
rect 380 -3180 640 -3140
<< viali >>
rect 1140 -20 1200 120
rect 380 -180 640 -140
rect 380 -300 640 -260
rect 1140 -620 1200 -480
rect 380 -780 640 -740
rect 380 -900 640 -860
rect 1140 -1220 1200 -1080
rect 380 -1380 640 -1340
rect 380 -1500 640 -1460
rect 1140 -1820 1200 -1680
rect 380 -1980 640 -1940
rect 380 -2100 640 -2060
rect 1140 -2420 1200 -2280
rect 380 -2580 640 -2540
rect 380 -2700 640 -2660
rect 1140 -3020 1200 -2880
rect 380 -3180 640 -3140
rect 380 -3300 640 -3260
rect 1140 -3620 1200 -3480
rect 380 -3780 640 -3740
rect 380 -3900 640 -3860
rect 1140 -4220 1200 -4080
rect 380 -4380 640 -4340
<< metal1 >>
rect 0 600 1400 800
rect 0 240 200 400
rect 0 180 1080 240
rect 0 0 200 180
rect 1140 140 1400 600
rect 380 120 480 140
rect 380 -40 400 120
rect 460 -40 480 120
rect 540 120 980 140
rect 540 -20 900 120
rect 960 -20 980 120
rect 540 -40 980 -20
rect 1040 120 1400 140
rect 1040 -20 1140 120
rect 1200 -20 1400 120
rect 380 -60 480 -40
rect 1040 -60 1400 -20
rect 300 -140 700 -120
rect 300 -180 380 -140
rect 640 -180 700 -140
rect 0 -360 200 -200
rect 300 -260 700 -180
rect 300 -300 380 -260
rect 640 -300 700 -260
rect 300 -320 700 -300
rect 0 -420 1080 -360
rect 0 -600 200 -420
rect 1140 -460 1400 -60
rect 380 -480 480 -460
rect 380 -640 400 -480
rect 460 -640 480 -480
rect 380 -660 480 -640
rect 540 -480 640 -460
rect 540 -640 560 -480
rect 620 -640 640 -480
rect 880 -480 980 -460
rect 880 -620 900 -480
rect 960 -620 980 -480
rect 880 -640 980 -620
rect 1040 -480 1400 -460
rect 1040 -620 1140 -480
rect 1200 -620 1400 -480
rect 540 -660 640 -640
rect 1040 -660 1400 -620
rect 300 -740 700 -720
rect 300 -780 380 -740
rect 640 -780 700 -740
rect 0 -960 200 -800
rect 300 -860 700 -780
rect 300 -900 380 -860
rect 640 -900 700 -860
rect 300 -920 700 -900
rect 0 -1020 1080 -960
rect 0 -1200 200 -1020
rect 1140 -1060 1400 -660
rect 380 -1080 480 -1060
rect 380 -1240 400 -1080
rect 460 -1240 480 -1080
rect 380 -1260 480 -1240
rect 540 -1080 640 -1060
rect 540 -1240 560 -1080
rect 620 -1240 640 -1080
rect 880 -1080 980 -1060
rect 880 -1220 900 -1080
rect 960 -1220 980 -1080
rect 880 -1240 980 -1220
rect 1040 -1080 1400 -1060
rect 1040 -1220 1140 -1080
rect 1200 -1220 1400 -1080
rect 540 -1260 640 -1240
rect 1040 -1260 1400 -1220
rect 300 -1340 700 -1320
rect 300 -1380 380 -1340
rect 640 -1380 700 -1340
rect 0 -1560 200 -1400
rect 300 -1460 700 -1380
rect 300 -1500 380 -1460
rect 640 -1500 700 -1460
rect 300 -1520 700 -1500
rect 0 -1620 1080 -1560
rect 0 -1800 200 -1620
rect 1140 -1660 1400 -1260
rect 380 -1680 480 -1660
rect 380 -1840 400 -1680
rect 460 -1840 480 -1680
rect 380 -1860 480 -1840
rect 540 -1680 640 -1660
rect 540 -1840 560 -1680
rect 620 -1840 640 -1680
rect 880 -1680 980 -1660
rect 880 -1820 900 -1680
rect 960 -1820 980 -1680
rect 880 -1840 980 -1820
rect 1040 -1680 1400 -1660
rect 1040 -1820 1140 -1680
rect 1200 -1820 1400 -1680
rect 540 -1860 640 -1840
rect 1040 -1860 1400 -1820
rect 300 -1940 700 -1920
rect 300 -1980 380 -1940
rect 640 -1980 700 -1940
rect 0 -2160 200 -2000
rect 300 -2060 700 -1980
rect 300 -2100 380 -2060
rect 640 -2100 700 -2060
rect 300 -2120 700 -2100
rect 0 -2220 1080 -2160
rect 0 -2400 200 -2220
rect 1140 -2260 1400 -1860
rect 1600 -1820 1800 -1800
rect 1600 -1980 1620 -1820
rect 1780 -1980 1800 -1820
rect 1600 -2000 1800 -1980
rect 380 -2280 480 -2260
rect 380 -2440 400 -2280
rect 460 -2440 480 -2280
rect 380 -2460 480 -2440
rect 540 -2280 640 -2260
rect 540 -2440 560 -2280
rect 620 -2440 640 -2280
rect 880 -2280 980 -2260
rect 880 -2420 900 -2280
rect 960 -2420 980 -2280
rect 880 -2440 980 -2420
rect 1040 -2280 1400 -2260
rect 1040 -2420 1140 -2280
rect 1200 -2420 1400 -2280
rect 540 -2460 640 -2440
rect 1040 -2460 1400 -2420
rect 300 -2540 700 -2520
rect 300 -2580 380 -2540
rect 640 -2580 700 -2540
rect 0 -2760 200 -2600
rect 300 -2660 700 -2580
rect 300 -2700 380 -2660
rect 640 -2700 700 -2660
rect 300 -2720 700 -2700
rect 0 -2820 1080 -2760
rect 0 -3000 200 -2820
rect 1140 -2860 1400 -2460
rect 380 -2880 480 -2860
rect 380 -3040 400 -2880
rect 460 -3040 480 -2880
rect 380 -3060 480 -3040
rect 540 -2880 640 -2860
rect 540 -3040 560 -2880
rect 620 -3040 640 -2880
rect 880 -2880 980 -2860
rect 880 -3020 900 -2880
rect 960 -3020 980 -2880
rect 880 -3040 980 -3020
rect 1040 -2880 1400 -2860
rect 1040 -3020 1140 -2880
rect 1200 -3020 1400 -2880
rect 540 -3060 640 -3040
rect 1040 -3060 1400 -3020
rect 300 -3140 700 -3120
rect 300 -3180 380 -3140
rect 640 -3180 700 -3140
rect 0 -3360 200 -3200
rect 300 -3260 700 -3180
rect 300 -3300 380 -3260
rect 640 -3300 700 -3260
rect 300 -3320 700 -3300
rect 0 -3420 1080 -3360
rect 0 -3600 200 -3420
rect 1140 -3460 1400 -3060
rect 380 -3480 480 -3460
rect 380 -3640 400 -3480
rect 460 -3640 480 -3480
rect 380 -3660 480 -3640
rect 540 -3480 640 -3460
rect 540 -3640 560 -3480
rect 620 -3640 640 -3480
rect 880 -3480 980 -3460
rect 880 -3620 900 -3480
rect 960 -3620 980 -3480
rect 880 -3640 980 -3620
rect 1040 -3480 1400 -3460
rect 1040 -3620 1140 -3480
rect 1200 -3620 1400 -3480
rect 540 -3660 640 -3640
rect 1040 -3660 1400 -3620
rect 300 -3740 700 -3720
rect 300 -3780 380 -3740
rect 640 -3780 700 -3740
rect 0 -3960 200 -3800
rect 300 -3860 700 -3780
rect 300 -3900 380 -3860
rect 640 -3900 700 -3860
rect 300 -3920 700 -3900
rect 0 -4020 1080 -3960
rect 0 -4200 200 -4020
rect 1140 -4060 1400 -3660
rect 380 -4082 480 -4060
rect 380 -4236 396 -4082
rect 468 -4236 480 -4082
rect 380 -4260 480 -4236
rect 540 -4320 700 -4060
rect 880 -4080 980 -4060
rect 880 -4220 900 -4080
rect 960 -4220 980 -4080
rect 880 -4240 980 -4220
rect 1040 -4080 1400 -4060
rect 1040 -4220 1140 -4080
rect 1200 -4220 1400 -4080
rect 1040 -4260 1400 -4220
rect 1140 -4300 1400 -4260
rect 300 -4340 700 -4320
rect 300 -4380 380 -4340
rect 640 -4380 700 -4340
rect 300 -4400 700 -4380
rect 0 -4600 700 -4400
<< via1 >>
rect 400 -40 460 120
rect 900 -20 960 120
rect 400 -640 460 -480
rect 560 -640 620 -480
rect 900 -620 960 -480
rect 400 -1240 460 -1080
rect 560 -1240 620 -1080
rect 900 -1220 960 -1080
rect 400 -1840 460 -1680
rect 560 -1840 620 -1680
rect 900 -1820 960 -1680
rect 1620 -1980 1780 -1820
rect 400 -2440 460 -2280
rect 560 -2440 620 -2280
rect 900 -2420 960 -2280
rect 400 -3040 460 -2880
rect 560 -3040 620 -2880
rect 900 -3020 960 -2880
rect 400 -3640 460 -3480
rect 560 -3640 620 -3480
rect 900 -3620 960 -3480
rect 396 -4236 468 -4082
rect 900 -4220 960 -4080
<< metal2 >>
rect 380 120 480 140
rect 380 -40 400 120
rect 460 -40 480 120
rect 380 -480 480 -40
rect 880 120 980 140
rect 880 -20 900 120
rect 960 -20 980 120
rect 380 -640 400 -480
rect 460 -640 480 -480
rect 380 -660 480 -640
rect 540 -480 640 -460
rect 540 -640 560 -480
rect 620 -640 640 -480
rect 380 -1080 480 -1060
rect 380 -1240 400 -1080
rect 460 -1240 480 -1080
rect 380 -1680 480 -1240
rect 540 -1080 640 -640
rect 540 -1240 560 -1080
rect 620 -1240 640 -1080
rect 540 -1260 640 -1240
rect 880 -480 980 -20
rect 880 -620 900 -480
rect 960 -620 980 -480
rect 880 -1080 980 -620
rect 880 -1220 900 -1080
rect 960 -1220 980 -1080
rect 380 -1840 400 -1680
rect 460 -1840 480 -1680
rect 380 -1860 480 -1840
rect 540 -1680 640 -1660
rect 540 -1840 560 -1680
rect 620 -1840 640 -1680
rect 380 -2280 480 -2260
rect 380 -2440 400 -2280
rect 460 -2440 480 -2280
rect 380 -2880 480 -2440
rect 540 -2280 640 -1840
rect 540 -2440 560 -2280
rect 620 -2440 640 -2280
rect 540 -2460 640 -2440
rect 880 -1680 980 -1220
rect 880 -1820 900 -1680
rect 960 -1800 980 -1680
rect 960 -1820 1800 -1800
rect 880 -1980 1620 -1820
rect 1780 -1980 1800 -1820
rect 880 -2000 1800 -1980
rect 880 -2280 980 -2000
rect 880 -2420 900 -2280
rect 960 -2420 980 -2280
rect 380 -3040 400 -2880
rect 460 -3040 480 -2880
rect 380 -3060 480 -3040
rect 540 -2880 640 -2860
rect 540 -3040 560 -2880
rect 620 -3040 640 -2880
rect 380 -3480 480 -3460
rect 380 -3640 400 -3480
rect 460 -3640 480 -3480
rect 380 -4082 480 -3640
rect 540 -3480 640 -3040
rect 540 -3640 560 -3480
rect 620 -3640 640 -3480
rect 540 -3660 640 -3640
rect 880 -2880 980 -2420
rect 880 -3020 900 -2880
rect 960 -3020 980 -2880
rect 880 -3480 980 -3020
rect 880 -3620 900 -3480
rect 960 -3620 980 -3480
rect 380 -4236 396 -4082
rect 468 -4236 480 -4082
rect 380 -4260 480 -4236
rect 880 -4080 980 -3620
rect 880 -4220 900 -4080
rect 960 -4220 980 -4080
rect 880 -4240 980 -4220
use sky130_fd_pr__nfet_01v8_64Z3AY  sky130_fd_pr__nfet_01v8_64Z3AY_0 ~/tt_analog_z2a_2/mag
timestamp 1769862601
transform 1 0 511 0 1 79
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  sky130_fd_pr__pfet_01v8_MGS3BN_0
timestamp 1769202985
transform 1 0 1011 0 1 -516
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM0
timestamp 1769862601
transform 1 0 511 0 1 -4121
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64Z3AY  XM1
timestamp 1769862601
transform 1 0 511 0 1 -3521
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64Z3AY  XM2
timestamp 1769862601
transform 1 0 511 0 1 -2921
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64Z3AY  XM3
timestamp 1769862601
transform 1 0 511 0 1 -2321
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64Z3AY  XM4
timestamp 1769862601
transform 1 0 511 0 1 -1721
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64Z3AY  XM5
timestamp 1769862601
transform 1 0 511 0 1 -1121
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64Z3AY  XM6
timestamp 1769862601
transform 1 0 511 0 1 -521
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM8
timestamp 1769202985
transform 1 0 1011 0 1 84
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_MGS3BN  XM10
timestamp 1769202985
transform 1 0 1011 0 1 -1116
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_MGS3BN  XM11
timestamp 1769202985
transform 1 0 1011 0 1 -1716
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_MGS3BN  XM12
timestamp 1769202985
transform 1 0 1011 0 1 -2316
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_MGS3BN  XM13
timestamp 1769202985
transform 1 0 1011 0 1 -2916
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_MGS3BN  XM14
timestamp 1769202985
transform 1 0 1011 0 1 -3516
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_MGS3BN  XM15
timestamp 1769202985
transform 1 0 1011 0 1 -4116
box -211 -284 211 284
<< labels >>
flabel metal1 0 -4100 200 -3900 0 FreeSans 256 0 0 0 NAND_IN_0
port 10 nsew
flabel metal1 0 -3500 200 -3300 0 FreeSans 256 0 0 0 NAND_IN_1
port 9 nsew
flabel metal1 0 100 200 300 0 FreeSans 256 0 0 0 NAND_IN_7
port 1 nsew
flabel metal1 0 -500 200 -300 0 FreeSans 256 0 0 0 NAND_IN_6
port 3 nsew
flabel metal1 0 -4600 200 -4400 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 0 -1100 200 -900 0 FreeSans 256 0 0 0 NAND_IN_5
port 5 nsew
flabel metal1 0 -1700 200 -1500 0 FreeSans 256 0 0 0 NAND_IN_4
port 6 nsew
flabel metal1 0 -2300 200 -2100 0 FreeSans 256 0 0 0 NAND_IN_3
port 7 nsew
flabel metal1 0 -2900 200 -2700 0 FreeSans 256 0 0 0 NAND_IN_2
port 8 nsew
flabel metal1 0 600 200 800 0 FreeSans 256 0 0 0 VDD
port 2 nsew
flabel metal1 1600 -2000 1800 -1800 0 FreeSans 256 0 0 0 NAND_OUT
port 0 nsew
<< end >>
