magic
tech sky130A
magscale 1 2
timestamp 1769863106
<< error_s >>
rect 6440 -1640 6449 -1631
rect 6771 -1640 6780 -1631
rect 6431 -1645 6789 -1640
rect 6431 -1649 6445 -1645
rect 6440 -2551 6445 -1649
rect 6431 -2555 6445 -2551
rect 6775 -1649 6789 -1645
rect 6775 -2551 6780 -1649
rect 6775 -2555 6789 -2551
rect 6431 -2560 6789 -2555
rect 6440 -2569 6449 -2560
rect 6771 -2569 6780 -2560
<< metal1 >>
rect 800 1800 5400 2000
rect 800 -1000 1000 1800
rect 4800 400 5200 600
rect 6400 400 6800 600
rect 1800 200 3400 400
rect 1800 -400 2000 200
rect 3200 -400 3400 -200
rect 6400 -260 6600 -200
rect 6040 -320 6600 -260
rect 1800 -800 2000 -600
rect 2600 -1200 3400 -800
rect 4600 -1200 5800 -800
rect 3000 -1800 3400 -1600
rect 6400 -1640 6600 -320
rect 800 -3800 1000 -3200
rect 1800 -3400 2000 -3000
rect 3000 -3400 3200 -1800
rect 4800 -2600 5200 -2400
rect 6400 -2560 6440 -1640
rect 6780 -2560 6800 -2400
rect 6400 -2600 6800 -2560
rect 1800 -3600 3200 -3400
rect 800 -4000 3400 -3800
rect 4000 -4000 6000 -3800
<< via1 >>
rect 3460 -380 3620 -220
rect 3420 -2380 3580 -2220
rect 6440 -2560 6780 -1640
<< metal2 >>
rect 3400 -220 3640 -200
rect 3400 -380 3460 -220
rect 3620 -380 3640 -220
rect 3400 -400 3640 -380
rect 3400 -2220 3600 -400
rect 6400 -1000 6600 600
rect 5400 -1200 6600 -1000
rect 5400 -1800 5600 -1200
rect 3400 -2380 3420 -2220
rect 3580 -2380 3600 -2220
rect 3400 -2400 3600 -2380
<< via2 >>
rect 6440 -2560 6780 -1640
use NAND2  x1
timestamp 1769862601
transform 1 0 3600 0 -1 -2200
box -200 -1200 1200 1800
use NAND2  x2
timestamp 1769862601
transform 1 0 5200 0 -1 -2200
box -200 -1200 1200 1800
use NAND2  x3
timestamp 1769862601
transform 1 0 3600 0 1 200
box -200 -1200 1200 1800
use NAND2  x4
timestamp 1769862601
transform 1 0 5200 0 1 200
box -200 -1200 1200 1800
use inv_x4  x24 ~/tt_analog_z2a_2/mag
timestamp 1769635883
transform 0 -1 1600 -1 0 400
box 800 -1200 3600 800
<< labels >>
flabel metal1 3200 -1200 3400 -1000 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 3200 1800 3400 2000 0 FreeSans 256 0 0 0 VDD
port 4 nsew
flabel metal1 3200 200 3400 400 0 FreeSans 256 0 0 0 T_IN
port 1 nsew
flabel metal1 3200 -400 3400 -200 0 FreeSans 256 0 0 0 CLK
port 2 nsew
flabel metal1 6400 400 6600 600 0 FreeSans 256 0 0 0 Q
port 0 nsew
flabel metal1 6400 -2600 6600 -2400 0 FreeSans 256 0 0 0 ZQ
port 3 nsew
<< end >>
