magic
tech sky130A
timestamp 1770560933
<< metal1 >>
rect 200 -2900 3900 -2800
rect 200 -3300 300 -3200
rect 600 -3210 700 -3200
rect 600 -3290 610 -3210
rect 690 -3290 700 -3210
rect 600 -3300 700 -3290
rect 800 -3210 900 -3200
rect 800 -3290 810 -3210
rect 890 -3290 900 -3210
rect 800 -3300 900 -3290
rect 1100 -3210 1200 -3200
rect 1100 -3290 1110 -3210
rect 1190 -3290 1200 -3210
rect 1100 -3300 1200 -3290
rect 1300 -3210 1400 -3200
rect 1300 -3290 1310 -3210
rect 1390 -3290 1400 -3210
rect 1300 -3300 1400 -3290
rect 1600 -3210 1700 -3200
rect 1600 -3290 1610 -3210
rect 1690 -3290 1700 -3210
rect 1600 -3300 1700 -3290
rect 1800 -3210 1900 -3200
rect 1800 -3290 1810 -3210
rect 1890 -3290 1900 -3210
rect 1800 -3300 1900 -3290
rect 2100 -3210 2200 -3200
rect 2100 -3290 2110 -3210
rect 2190 -3290 2200 -3210
rect 2100 -3300 2200 -3290
rect 2300 -3210 2400 -3200
rect 2300 -3290 2310 -3210
rect 2390 -3290 2400 -3210
rect 2300 -3300 2400 -3290
rect 2600 -3210 2700 -3200
rect 2600 -3290 2610 -3210
rect 2690 -3290 2700 -3210
rect 2600 -3300 2700 -3290
rect 2800 -3210 2900 -3200
rect 2800 -3290 2810 -3210
rect 2890 -3290 2900 -3210
rect 2800 -3300 2900 -3290
rect 3100 -3210 3200 -3200
rect 3100 -3290 3110 -3210
rect 3190 -3290 3200 -3210
rect 3100 -3300 3200 -3290
rect 3400 -3300 3500 -3200
rect 3600 -3210 3700 -3200
rect 3600 -3290 3610 -3210
rect 3690 -3290 3700 -3210
rect 3600 -3300 3700 -3290
rect 3800 -3210 3900 -3200
rect 3800 -3290 3810 -3210
rect 3890 -3290 3900 -3210
rect 3800 -3300 3900 -3290
rect 4200 -3210 4300 -3200
rect 4200 -3290 4210 -3210
rect 4290 -3290 4300 -3210
rect 4200 -3300 4300 -3290
rect 200 -3700 300 -3600
rect 400 -3700 800 -3600
rect 900 -3700 1300 -3600
rect 1400 -3700 1800 -3600
rect 1900 -3700 2300 -3600
rect 2400 -3700 2800 -3600
rect 2900 -3700 3300 -3600
rect 3400 -3700 3800 -3600
rect 600 -3810 700 -3800
rect 600 -3890 610 -3810
rect 690 -3890 700 -3810
rect 600 -3900 700 -3890
rect 1100 -3810 1200 -3800
rect 1100 -3890 1110 -3810
rect 1190 -3890 1200 -3810
rect -200 -4710 -150 -4700
rect -200 -4740 -190 -4710
rect -160 -4740 -150 -4710
rect -200 -4850 -150 -4740
rect -100 -4710 -50 -4700
rect -100 -4740 -90 -4710
rect -60 -4740 -50 -4710
rect -100 -4850 -50 -4740
rect 0 -4710 50 -4700
rect 0 -4740 10 -4710
rect 40 -4740 50 -4710
rect 0 -4850 50 -4740
rect 100 -4710 150 -4700
rect 100 -4740 110 -4710
rect 140 -4740 150 -4710
rect 100 -4850 150 -4740
rect 200 -4710 250 -4700
rect 200 -4740 210 -4710
rect 240 -4740 250 -4710
rect 200 -4850 250 -4740
rect 300 -4710 350 -4700
rect 300 -4740 310 -4710
rect 340 -4740 350 -4710
rect 300 -4850 350 -4740
rect 400 -4710 450 -4700
rect 400 -4740 410 -4710
rect 440 -4740 450 -4710
rect 400 -4850 450 -4740
rect 500 -4710 550 -4700
rect 500 -4740 510 -4710
rect 540 -4740 550 -4710
rect 500 -4850 550 -4740
rect 600 -4750 650 -3900
rect 1100 -3950 1200 -3890
rect 700 -4000 1200 -3950
rect 1600 -3810 1700 -3800
rect 1600 -3890 1610 -3810
rect 1690 -3890 1700 -3810
rect 700 -4750 750 -4000
rect 1600 -4050 1700 -3890
rect 800 -4100 1700 -4050
rect 2100 -3810 2200 -3800
rect 2100 -3890 2110 -3810
rect 2190 -3890 2200 -3810
rect 800 -4750 850 -4100
rect 2100 -4150 2200 -3890
rect 900 -4200 2200 -4150
rect 2600 -3810 2700 -3800
rect 2600 -3890 2610 -3810
rect 2690 -3890 2700 -3810
rect 900 -4750 950 -4200
rect 2600 -4250 2700 -3890
rect 1000 -4300 2700 -4250
rect 3100 -3810 3200 -3800
rect 3100 -3890 3110 -3810
rect 3190 -3890 3200 -3810
rect 3100 -4300 3200 -3890
rect 1000 -4750 1050 -4300
rect 2900 -4350 3200 -4300
rect 1100 -4400 3200 -4350
rect 3600 -3810 3700 -3800
rect 3600 -3890 3610 -3810
rect 3690 -3890 3700 -3810
rect 3600 -4400 3700 -3890
rect 1100 -4750 1150 -4400
rect 3400 -4450 3700 -4400
rect 1200 -4500 3700 -4450
rect 4200 -3810 4300 -3800
rect 4200 -3890 4210 -3810
rect 4290 -3890 4300 -3810
rect 1200 -4750 1250 -4500
rect 4200 -4550 4300 -3890
rect 1300 -4600 4300 -4550
rect 1300 -4750 1350 -4600
<< via1 >>
rect 310 -3290 390 -3210
rect 610 -3290 690 -3210
rect 810 -3290 890 -3210
rect 1110 -3290 1190 -3210
rect 1310 -3290 1390 -3210
rect 1610 -3290 1690 -3210
rect 1810 -3290 1890 -3210
rect 2110 -3290 2190 -3210
rect 2310 -3290 2390 -3210
rect 2610 -3290 2690 -3210
rect 2810 -3290 2890 -3210
rect 3110 -3290 3190 -3210
rect 3310 -3290 3390 -3210
rect 3610 -3290 3690 -3210
rect 3810 -3290 3890 -3210
rect 4210 -3290 4290 -3210
rect 610 -3890 690 -3810
rect 1110 -3890 1190 -3810
rect -190 -4740 -160 -4710
rect -90 -4740 -60 -4710
rect 10 -4740 40 -4710
rect 110 -4740 140 -4710
rect 210 -4740 240 -4710
rect 310 -4740 340 -4710
rect 410 -4740 440 -4710
rect 510 -4740 540 -4710
rect 1610 -3890 1690 -3810
rect 2110 -3890 2190 -3810
rect 2610 -3890 2690 -3810
rect 3110 -3890 3190 -3810
rect 3610 -3890 3690 -3810
rect 4210 -3890 4290 -3810
<< metal2 >>
rect 300 -3210 400 -2700
rect 300 -3290 310 -3210
rect 390 -3290 400 -3210
rect 300 -3850 400 -3290
rect -200 -3900 400 -3850
rect 600 -3210 700 -3200
rect 600 -3290 610 -3210
rect 690 -3290 700 -3210
rect 600 -3810 700 -3290
rect 600 -3890 610 -3810
rect 690 -3890 700 -3810
rect 600 -3900 700 -3890
rect 800 -3210 900 -2700
rect 800 -3290 810 -3210
rect 890 -3290 900 -3210
rect -200 -4710 -150 -3900
rect 800 -3950 900 -3290
rect 1100 -3210 1200 -3200
rect 1100 -3290 1110 -3210
rect 1190 -3290 1200 -3210
rect 1100 -3810 1200 -3290
rect 1100 -3890 1110 -3810
rect 1190 -3890 1200 -3810
rect 1100 -3900 1200 -3890
rect 1300 -3210 1400 -2700
rect 1300 -3290 1310 -3210
rect 1390 -3290 1400 -3210
rect -200 -4740 -190 -4710
rect -160 -4740 -150 -4710
rect -200 -4750 -150 -4740
rect -100 -4000 900 -3950
rect -100 -4710 -50 -4000
rect 1300 -4050 1400 -3290
rect 1600 -3210 1700 -3200
rect 1600 -3290 1610 -3210
rect 1690 -3290 1700 -3210
rect 1600 -3810 1700 -3290
rect 1600 -3890 1610 -3810
rect 1690 -3890 1700 -3810
rect 1600 -3900 1700 -3890
rect 1800 -3210 1900 -2700
rect 1800 -3290 1810 -3210
rect 1890 -3290 1900 -3210
rect -100 -4740 -90 -4710
rect -60 -4740 -50 -4710
rect -100 -4750 -50 -4740
rect 0 -4100 1400 -4050
rect 0 -4710 50 -4100
rect 1800 -4150 1900 -3290
rect 2100 -3210 2200 -3200
rect 2100 -3290 2110 -3210
rect 2190 -3290 2200 -3210
rect 2100 -3810 2200 -3290
rect 2100 -3890 2110 -3810
rect 2190 -3890 2200 -3810
rect 2100 -3900 2200 -3890
rect 2300 -3210 2400 -2700
rect 2300 -3290 2310 -3210
rect 2390 -3290 2400 -3210
rect 0 -4740 10 -4710
rect 40 -4740 50 -4710
rect 0 -4750 50 -4740
rect 100 -4200 1900 -4150
rect 100 -4710 150 -4200
rect 2300 -4250 2400 -3290
rect 2600 -3210 2700 -3200
rect 2600 -3290 2610 -3210
rect 2690 -3290 2700 -3210
rect 2600 -3810 2700 -3290
rect 2600 -3890 2610 -3810
rect 2690 -3890 2700 -3810
rect 2600 -3900 2700 -3890
rect 2800 -3210 2900 -2700
rect 2800 -3290 2810 -3210
rect 2890 -3290 2900 -3210
rect 100 -4740 110 -4710
rect 140 -4740 150 -4710
rect 100 -4750 150 -4740
rect 200 -4300 2400 -4250
rect 200 -4710 250 -4300
rect 2800 -4350 2900 -3290
rect 3100 -3210 3200 -3200
rect 3100 -3290 3110 -3210
rect 3190 -3290 3200 -3210
rect 3100 -3810 3200 -3290
rect 3100 -3890 3110 -3810
rect 3190 -3890 3200 -3810
rect 3100 -3900 3200 -3890
rect 3300 -3210 3400 -2700
rect 3300 -3290 3310 -3210
rect 3390 -3290 3400 -3210
rect 200 -4740 210 -4710
rect 240 -4740 250 -4710
rect 200 -4750 250 -4740
rect 300 -4400 2900 -4350
rect 300 -4710 350 -4400
rect 3300 -4450 3400 -3290
rect 3600 -3210 3700 -3200
rect 3600 -3290 3610 -3210
rect 3690 -3290 3700 -3210
rect 3600 -3810 3700 -3290
rect 3600 -3890 3610 -3810
rect 3690 -3890 3700 -3810
rect 3600 -3900 3700 -3890
rect 3800 -3210 3900 -2700
rect 3800 -3290 3810 -3210
rect 3890 -3290 3900 -3210
rect 300 -4740 310 -4710
rect 340 -4740 350 -4710
rect 300 -4750 350 -4740
rect 400 -4500 3400 -4450
rect 400 -4710 450 -4500
rect 3800 -4550 3900 -3290
rect 4200 -3210 4300 -3200
rect 4200 -3290 4210 -3210
rect 4290 -3290 4300 -3210
rect 4200 -3810 4300 -3290
rect 4200 -3890 4210 -3810
rect 4290 -3890 4300 -3810
rect 4200 -3900 4300 -3890
rect 400 -4740 410 -4710
rect 440 -4740 450 -4710
rect 400 -4750 450 -4740
rect 500 -4600 3900 -4550
rect 500 -4710 550 -4600
rect 500 -4740 510 -4710
rect 540 -4740 550 -4710
rect 500 -4750 550 -4740
use inv_x1  x1 ~/tt_analog_z2a_2/mag
timestamp 1770560933
transform 1 0 200 0 1 -3000
box 100 -700 500 200
use inv_x1  x2
timestamp 1770560933
transform 1 0 700 0 1 -3000
box 100 -700 500 200
use inv_x1  x3
timestamp 1770560933
transform 1 0 1200 0 1 -3000
box 100 -700 500 200
use inv_x1  x4
timestamp 1770560933
transform 1 0 1700 0 1 -3000
box 100 -700 500 200
use inv_x1  x5
timestamp 1770560933
transform 1 0 2200 0 1 -3000
box 100 -700 500 200
use inv_x1  x6
timestamp 1770560933
transform 1 0 2700 0 1 -3000
box 100 -700 500 200
use inv_x1  x7
timestamp 1770560933
transform 1 0 3200 0 1 -3000
box 100 -700 500 200
use inv_x1  x28
timestamp 1770560933
transform 1 0 3700 0 1 -3000
box 100 -700 500 200
<< labels >>
flabel metal1 200 -3700 300 -3600 0 FreeSans 128 0 0 0 VSS
port 18 nsew
flabel metal1 200 -2900 300 -2800 0 FreeSans 128 0 0 0 VDD
port 17 nsew
flabel metal1 200 -3300 300 -3200 0 FreeSans 128 0 0 0 LOGICIN_0_2
port 15 nsew
flabel metal1 600 -3300 700 -3200 0 FreeSans 128 0 0 0 Z_LOGICIN_0_2
port 16 nsew
flabel metal1 1100 -3300 1200 -3200 0 FreeSans 128 0 0 0 Z_LOGICIN_0_4
port 14 nsew
flabel metal1 800 -3300 900 -3200 0 FreeSans 128 0 0 0 LOGICIN_0_4
port 13 nsew
flabel metal1 1300 -3300 1400 -3200 0 FreeSans 128 0 0 0 LOGICIN_0_6
port 12 nsew
flabel metal1 3800 -3300 3900 -3200 0 FreeSans 128 0 0 0 LOGICIN_1_6
port 0 nsew
flabel metal1 3600 -3300 3700 -3200 0 FreeSans 128 0 0 0 Z_LOGICIN_1_4
port 2 nsew
flabel metal1 3400 -3300 3500 -3200 0 FreeSans 128 0 0 0 LOGICIN_1_4
port 3 nsew
flabel metal1 2800 -3300 2900 -3200 0 FreeSans 128 0 0 0 LOGICIN_1_2
port 4 nsew
flabel metal1 3100 -3300 3200 -3200 0 FreeSans 128 0 0 0 Z_LOGICIN_1_2
port 5 nsew
flabel metal1 2300 -3300 2400 -3200 0 FreeSans 128 0 0 0 LOGICIN_1_0
port 6 nsew
flabel metal1 2600 -3300 2700 -3200 0 FreeSans 128 0 0 0 Z_LOGICIN_1_0
port 7 nsew
flabel metal1 2100 -3300 2200 -3200 0 FreeSans 128 0 0 0 Z_LOGICIN_0_8
port 9 nsew
flabel metal1 1600 -3300 1700 -3200 0 FreeSans 128 0 0 0 Z_LOGICIN_0_6
port 11 nsew
flabel metal1 1800 -3300 1900 -3200 0 FreeSans 128 0 0 0 LOGICIN_0_8
port 10 nsew
flabel metal1 4200 -3300 4300 -3200 0 FreeSans 128 0 0 0 Z_LOGICIN_1_6
port 1 nsew
<< end >>
