magic
tech sky130A
timestamp 1770560933
<< metal1 >>
rect 300 300 400 400
rect -100 50 200 100
rect -100 -150 -50 50
rect 150 0 200 50
rect 7200 50 7500 100
rect 150 -100 300 0
rect 150 -150 200 -100
rect -100 -200 200 -150
rect 7200 -150 7250 50
rect 7450 -150 7500 50
rect 7200 -200 7500 -150
rect 300 -400 400 -300
<< via1 >>
rect -50 -150 150 50
rect 7250 -150 7450 50
<< metal2 >>
rect -100 50 7500 100
rect -100 -150 -50 50
rect 150 -150 7250 50
rect 7450 -150 7500 50
rect -100 -200 7500 -150
use inv_x4  x7 ~/tt_analog_z2a_2/mag
timestamp 1770560933
transform 1 0 -100 0 1 100
box 400 -600 1800 400
use inv_x4  x9
timestamp 1770560933
transform 1 0 1300 0 1 100
box 400 -600 1800 400
use inv_x4  x10
timestamp 1770560933
transform 1 0 2700 0 1 100
box 400 -600 1800 400
use inv_x4  x11
timestamp 1770560933
transform 1 0 4100 0 1 100
box 400 -600 1800 400
use inv_x4  x12
timestamp 1770560933
transform 1 0 5500 0 1 100
box 400 -600 1800 400
<< labels >>
flabel metal1 300 300 400 400 0 FreeSans 128 0 0 0 VDD
port 0 nsew
flabel metal1 300 -400 400 -300 0 FreeSans 128 0 0 0 VSS
port 1 nsew
flabel via1 7300 -100 7400 0 0 FreeSans 128 0 0 0 OUT_OSC5
port 2 nsew
<< end >>
