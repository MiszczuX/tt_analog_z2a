magic
tech sky130A
magscale 1 2
timestamp 1769198914
<< metal1 >>
rect -5800 3400 -1400 3600
rect -5800 -700 -5000 3400
rect -2800 2600 -1600 2800
rect 6200 1800 8000 2000
rect -2900 1300 -2700 1400
rect -2900 1280 -2000 1300
rect -2900 1220 -2180 1280
rect -2020 1220 -2000 1280
rect -2900 1200 -2000 1220
rect -3200 1100 -3000 1200
rect -3200 1080 -1800 1100
rect -3200 1020 -1980 1080
rect -1820 1020 -1800 1080
rect -3200 1000 -1800 1020
rect -3500 900 -3300 1000
rect -3500 880 -1600 900
rect -3500 820 -1780 880
rect -1620 820 -1600 880
rect -3500 800 -1600 820
rect -3800 700 -3600 800
rect -3800 680 -1400 700
rect -3800 620 -1580 680
rect -1420 620 -1400 680
rect -3800 600 -1400 620
rect -3600 480 -1200 500
rect -3600 420 -1380 480
rect -1220 420 -1200 480
rect -3600 400 -1200 420
rect -3600 300 -3400 400
rect -3300 280 -1000 300
rect -3300 220 -1180 280
rect -1020 220 -1000 280
rect -3300 200 -1000 220
rect 7800 200 8000 1800
rect -3300 100 -3100 200
rect -3000 80 -860 100
rect -3000 20 -980 80
rect -880 20 -860 80
rect -3000 0 -860 20
rect 7000 0 8000 200
rect -3000 -100 -2800 0
rect -5800 -2500 -5700 -700
rect -5100 -2500 -5000 -700
rect -3000 -800 -2600 -600
rect -3000 -1300 -2600 -1100
rect -3000 -1900 -2600 -1700
rect -3000 -2500 -2600 -2300
rect -5800 -2600 -5000 -2500
rect -3000 -3100 -2600 -2900
rect -3000 -3700 -2600 -3500
rect -3000 -4300 -2600 -4100
rect -3000 -4900 -2600 -4700
rect -3000 -5500 -2600 -5300
rect -2400 -5320 -2300 -500
rect -2400 -5480 -2380 -5320
rect -2320 -5480 -2300 -5320
rect -3000 -6200 -2600 -5800
rect -3000 -6700 -2600 -6500
rect -2400 -6540 -2300 -5480
rect -2400 -6680 -2380 -6540
rect -2320 -6680 -2300 -6540
rect -3000 -7300 -2600 -7100
rect -3000 -7900 -2600 -7700
rect -3000 -8500 -2600 -8300
rect -3000 -9100 -2600 -8900
rect -3000 -9700 -2600 -9500
rect -3000 -10300 -2600 -10100
rect -3000 -10900 -2600 -10700
rect -3000 -12100 -2600 -11900
rect -3000 -12700 -2600 -12500
rect -3000 -13300 -2600 -13100
rect -3000 -13900 -2600 -13700
rect -3000 -14500 -2600 -14300
rect -3000 -15100 -2600 -14900
rect -3000 -15700 -2600 -15500
rect -3000 -16300 -2600 -16100
rect -2400 -16120 -2300 -6680
rect -2400 -16280 -2380 -16120
rect -2320 -16280 -2300 -16120
rect -3000 -17500 -2600 -17300
rect -2400 -17320 -2300 -16280
rect -2400 -17480 -2380 -17320
rect -2320 -17480 -2300 -17320
rect -3000 -18100 -2600 -17900
rect -3000 -18700 -2600 -18500
rect -3000 -19300 -2600 -19100
rect -3000 -19900 -2600 -19700
rect -3000 -20500 -2600 -20300
rect -3000 -21100 -2600 -20900
rect -6788 -21804 -4192 -21542
rect -3000 -21700 -2600 -21500
rect -2400 -21800 -2300 -17480
rect -2200 -4720 -2100 -500
rect -2200 -4880 -2180 -4720
rect -2120 -4880 -2100 -4720
rect -2200 -7120 -2100 -4880
rect -2200 -7260 -2180 -7120
rect -2120 -7260 -2100 -7120
rect -2200 -15520 -2100 -7260
rect -2200 -15680 -2180 -15520
rect -2120 -15680 -2100 -15520
rect -2200 -17920 -2100 -15680
rect -2200 -18080 -2180 -17920
rect -2120 -18080 -2100 -17920
rect -2200 -21800 -2100 -18080
rect -2000 -4120 -1900 -500
rect -2000 -4280 -1980 -4120
rect -1920 -4280 -1900 -4120
rect -2000 -7720 -1900 -4280
rect -2000 -7880 -1980 -7720
rect -1920 -7880 -1900 -7720
rect -2000 -14920 -1900 -7880
rect -2000 -15080 -1980 -14920
rect -1920 -15080 -1900 -14920
rect -2000 -18520 -1900 -15080
rect -2000 -18680 -1980 -18520
rect -1920 -18680 -1900 -18520
rect -2000 -21800 -1900 -18680
rect -1800 -3520 -1700 -500
rect -1800 -3680 -1780 -3520
rect -1720 -3680 -1700 -3520
rect -1800 -8320 -1700 -3680
rect -1800 -8480 -1780 -8320
rect -1720 -8480 -1700 -8320
rect -1800 -14320 -1700 -8480
rect -1800 -14480 -1780 -14320
rect -1720 -14480 -1700 -14320
rect -1800 -19120 -1700 -14480
rect -1800 -19280 -1780 -19120
rect -1720 -19280 -1700 -19120
rect -1800 -21800 -1700 -19280
rect -1600 -2920 -1500 -500
rect -1600 -3080 -1580 -2920
rect -1520 -3080 -1500 -2920
rect -1600 -8920 -1500 -3080
rect -1600 -9080 -1580 -8920
rect -1520 -9080 -1500 -8920
rect -1600 -13720 -1500 -9080
rect -1600 -13880 -1580 -13720
rect -1520 -13880 -1500 -13720
rect -1600 -19720 -1500 -13880
rect -1600 -19880 -1580 -19720
rect -1520 -19880 -1500 -19720
rect -1600 -21800 -1500 -19880
rect -1400 -9520 -1300 -500
rect -1400 -9680 -1380 -9520
rect -1320 -9680 -1300 -9520
rect -1400 -13120 -1300 -9680
rect -1400 -13280 -1380 -13120
rect -1320 -13280 -1300 -13120
rect -1400 -20320 -1300 -13280
rect -1400 -20480 -1380 -20320
rect -1320 -20480 -1300 -20320
rect -1400 -21800 -1300 -20480
rect -1200 -12520 -1100 -500
rect -1200 -12680 -1180 -12520
rect -1120 -12680 -1100 -12520
rect -1200 -20920 -1100 -12680
rect -1200 -21080 -1180 -20920
rect -1120 -21080 -1100 -20920
rect -1200 -21800 -1100 -21080
rect -1000 -21520 -900 -500
rect -1000 -21680 -980 -21520
rect -920 -21680 -900 -21520
rect -1000 -21800 -900 -21680
rect -800 -21800 -700 -200
rect -600 -4720 -500 -300
rect -600 -4880 -580 -4720
rect -520 -4880 -500 -4720
rect -600 -21800 -500 -4880
rect -400 -4120 -300 -300
rect -400 -4280 -380 -4120
rect -320 -4280 -300 -4120
rect -400 -7720 -300 -4280
rect -400 -7880 -380 -7720
rect -320 -7880 -300 -7720
rect -400 -21800 -300 -7880
rect -200 -3520 -100 -300
rect -200 -3680 -180 -3520
rect -120 -3680 -100 -3520
rect -200 -8320 -100 -3680
rect -200 -8480 -180 -8320
rect -120 -8480 -100 -8320
rect -200 -14320 -100 -8480
rect -200 -14480 -180 -14320
rect -120 -14480 -100 -14320
rect -200 -21800 -100 -14480
rect 0 -2920 100 -300
rect 0 -3080 20 -2920
rect 80 -3080 100 -2920
rect 0 -8920 100 -3080
rect 0 -9080 20 -8920
rect 80 -9080 100 -8920
rect 0 -13720 100 -9080
rect 0 -13880 20 -13720
rect 80 -13880 100 -13720
rect 0 -17300 100 -13880
rect 200 -2320 300 -300
rect 200 -2480 220 -2320
rect 280 -2480 300 -2320
rect 200 -9520 300 -2480
rect 200 -9680 220 -9520
rect 280 -9680 300 -9520
rect 200 -13120 300 -9680
rect 200 -13280 220 -13120
rect 280 -13280 300 -13120
rect 0 -19720 100 -17500
rect 200 -17900 300 -13280
rect 400 -1720 500 -300
rect 400 -1880 420 -1720
rect 480 -1880 500 -1720
rect 400 -6500 500 -1880
rect 600 -1120 700 -300
rect 1000 -800 1200 -600
rect 3200 -800 3600 -600
rect 600 -1280 620 -1120
rect 680 -1280 700 -1120
rect 400 -6700 480 -6500
rect 400 -10120 500 -6700
rect 400 -10280 420 -10120
rect 480 -10280 500 -10120
rect 400 -12520 500 -10280
rect 400 -12680 420 -12520
rect 480 -12680 500 -12520
rect 0 -19880 20 -19720
rect 80 -19880 100 -19720
rect 0 -21800 100 -19880
rect 200 -20320 300 -18100
rect 200 -20480 220 -20320
rect 280 -20480 300 -20320
rect 200 -21800 300 -20480
rect 400 -20920 500 -12680
rect 400 -21080 420 -20920
rect 480 -21080 500 -20920
rect 400 -21800 500 -21080
rect 600 -10720 700 -1280
rect 3800 -3400 4000 -3200
rect 800 -4900 1000 -4800
rect 3600 -8000 3800 -4000
rect 6228 -5266 8358 -4896
rect 6228 -5602 6776 -5266
rect 7550 -5602 8358 -5266
rect 6228 -7464 8358 -5602
rect 4000 -8800 4200 -8600
rect 600 -10880 620 -10720
rect 680 -10880 700 -10720
rect 600 -11920 700 -10880
rect 600 -12080 620 -11920
rect 680 -12080 700 -11920
rect 600 -21520 700 -12080
rect 3800 -14200 4000 -14000
rect 1000 -17000 1200 -16800
rect 900 -17500 1000 -17300
rect 900 -18100 1100 -17900
rect 900 -18700 1100 -18500
rect 3600 -18800 3800 -14800
rect 900 -19300 1100 -19100
rect 3800 -19600 4000 -19400
rect 600 -21680 620 -21520
rect 680 -21680 700 -21520
rect 600 -21800 700 -21680
rect -6788 -22390 -6268 -21804
rect -4744 -21994 -4192 -21804
rect -4744 -22000 -2596 -21994
rect -4744 -22200 1200 -22000
rect -4744 -22390 -2596 -22200
rect -6788 -22474 -2596 -22390
rect -6788 -22720 -4192 -22474
<< via1 >>
rect -1380 2620 -1220 2780
rect -2180 1220 -2020 1280
rect -1980 1020 -1820 1080
rect -1780 820 -1620 880
rect -1580 620 -1420 680
rect -1380 420 -1220 480
rect -1180 220 -1020 280
rect 7000 200 7800 1800
rect -980 20 -880 80
rect -5700 -2500 -5100 -700
rect -2380 -5480 -2320 -5320
rect -2380 -6680 -2320 -6540
rect -2380 -16280 -2320 -16120
rect -2380 -17480 -2320 -17320
rect -2180 -4880 -2120 -4720
rect -2180 -7260 -2120 -7120
rect -2180 -15680 -2120 -15520
rect -2180 -18080 -2120 -17920
rect -1980 -4280 -1920 -4120
rect -1980 -7880 -1920 -7720
rect -1980 -15080 -1920 -14920
rect -1980 -18680 -1920 -18520
rect -1780 -3680 -1720 -3520
rect -1780 -8480 -1720 -8320
rect -1780 -14480 -1720 -14320
rect -1780 -19280 -1720 -19120
rect -1580 -3080 -1520 -2920
rect -1580 -9080 -1520 -8920
rect -1580 -13880 -1520 -13720
rect -1580 -19880 -1520 -19720
rect -1380 -9680 -1320 -9520
rect -1380 -13280 -1320 -13120
rect -1380 -20480 -1320 -20320
rect -1180 -12680 -1120 -12520
rect -1180 -21080 -1120 -20920
rect -980 -21680 -920 -21520
rect -580 -4880 -520 -4720
rect -380 -4280 -320 -4120
rect -380 -7880 -320 -7720
rect -180 -3680 -120 -3520
rect -180 -8480 -120 -8320
rect -180 -14480 -120 -14320
rect 20 -3080 80 -2920
rect 20 -9080 80 -8920
rect 20 -13880 80 -13720
rect 220 -2480 280 -2320
rect 220 -9680 280 -9520
rect 220 -13280 280 -13120
rect 420 -1880 480 -1720
rect 620 -1280 680 -1120
rect 420 -10280 480 -10120
rect 420 -12680 480 -12520
rect 20 -19880 80 -19720
rect 220 -20480 280 -20320
rect 420 -21080 480 -20920
rect 3200 -7800 3600 -4200
rect 6776 -5602 7550 -5266
rect 620 -10880 680 -10720
rect 620 -12080 680 -11920
rect 3200 -18600 3600 -15000
rect 620 -21680 680 -21520
rect -6268 -22390 -4744 -21804
<< metal2 >>
rect 6800 1800 8000 2000
rect 7800 200 8000 1800
rect -5544 -600 -2702 -520
rect -5800 -700 1200 -600
rect -5800 -1260 -5700 -700
rect -6494 -2500 -5700 -1260
rect -5100 -800 1200 -700
rect -5100 -970 -2702 -800
rect -5100 -1260 -5000 -970
rect -3400 -1120 1400 -1100
rect -5100 -2500 -4548 -1260
rect -3400 -1280 620 -1120
rect 680 -1280 1400 -1120
rect -3400 -1300 1400 -1280
rect -3400 -1720 1400 -1700
rect -3400 -1880 420 -1720
rect 480 -1880 1400 -1720
rect -3400 -1900 1400 -1880
rect -3400 -2320 1400 -2300
rect -3400 -2480 220 -2320
rect 280 -2480 1400 -2320
rect -3400 -2500 1400 -2480
rect -6494 -11106 -4548 -2500
rect -3400 -2920 -1500 -2900
rect -3400 -3080 -1580 -2920
rect -1520 -3080 -1500 -2920
rect -3400 -3100 -1500 -3080
rect 0 -2920 1400 -2900
rect 0 -3080 20 -2920
rect 80 -3080 1400 -2920
rect 0 -3100 1400 -3080
rect -3400 -3520 -1700 -3500
rect -3400 -3680 -1780 -3520
rect -1720 -3680 -1700 -3520
rect -3400 -3700 -1700 -3680
rect -200 -3520 1400 -3500
rect -200 -3680 -180 -3520
rect -120 -3680 1400 -3520
rect -200 -3700 1400 -3680
rect 7000 -4000 8000 200
rect -3400 -4120 -1900 -4100
rect -3400 -4280 -1980 -4120
rect -1920 -4280 -1900 -4120
rect -3400 -4300 -1900 -4280
rect -400 -4120 1400 -4100
rect -400 -4280 -380 -4120
rect -320 -4280 1400 -4120
rect -400 -4300 1400 -4280
rect 3000 -4200 8000 -4000
rect -3400 -4720 -2100 -4700
rect -3400 -4880 -2180 -4720
rect -2120 -4880 -2100 -4720
rect -3400 -4900 -2100 -4880
rect -600 -4720 1400 -4700
rect -600 -4880 -580 -4720
rect -520 -4880 1400 -4720
rect -600 -4900 1400 -4880
rect -3400 -5320 1400 -5300
rect -3400 -5480 -2380 -5320
rect -2320 -5480 1400 -5320
rect -3400 -5500 1400 -5480
rect -3000 -6200 1000 -5800
rect -3400 -6540 1400 -6500
rect -3400 -6680 -2380 -6540
rect -2320 -6680 1400 -6540
rect -3400 -6700 1400 -6680
rect -3400 -7120 1400 -7100
rect -3400 -7260 -2180 -7120
rect -2120 -7260 1400 -7120
rect -3400 -7300 1400 -7260
rect -3400 -7720 -1900 -7700
rect -3400 -7880 -1980 -7720
rect -1920 -7880 -1900 -7720
rect -3400 -7900 -1900 -7880
rect -400 -7720 1400 -7700
rect -400 -7880 -380 -7720
rect -320 -7880 1400 -7720
rect -400 -7900 1400 -7880
rect 3000 -7800 3200 -4200
rect 3600 -5266 8000 -4200
rect 3600 -5602 6776 -5266
rect 7550 -5602 8000 -5266
rect 3600 -6000 8000 -5602
rect 3600 -7800 3800 -6000
rect 3000 -8000 3800 -7800
rect -3400 -8320 -1700 -8300
rect -3400 -8480 -1780 -8320
rect -1720 -8480 -1700 -8320
rect -3400 -8500 -1700 -8480
rect -200 -8320 1400 -8300
rect -200 -8480 -180 -8320
rect -120 -8480 1400 -8320
rect -200 -8500 1400 -8480
rect -3400 -8920 -1500 -8900
rect -3400 -9080 -1580 -8920
rect -1520 -9080 -1500 -8920
rect -3400 -9100 -1500 -9080
rect 0 -8920 1400 -8900
rect 0 -9080 20 -8920
rect 80 -9080 1400 -8920
rect 0 -9100 1400 -9080
rect -3400 -9520 -1300 -9500
rect -3400 -9680 -1380 -9520
rect -1320 -9680 -1300 -9520
rect -3400 -9700 -1300 -9680
rect 200 -9520 1400 -9500
rect 200 -9680 220 -9520
rect 280 -9680 1400 -9520
rect 200 -9700 1400 -9680
rect -3400 -10120 1400 -10100
rect -3400 -10280 420 -10120
rect 480 -10280 1400 -10120
rect -3400 -10300 1400 -10280
rect -3400 -10720 1400 -10700
rect -3400 -10880 620 -10720
rect 680 -10880 1400 -10720
rect -3400 -10900 1400 -10880
rect -6494 -11200 -2914 -11106
rect -6494 -11600 1400 -11200
rect -6494 -11678 -2914 -11600
rect -6494 -21804 -4548 -11678
rect -3400 -11920 1400 -11900
rect -3400 -12080 620 -11920
rect 680 -12080 1400 -11920
rect -3400 -12100 1400 -12080
rect -3400 -12520 -1100 -12500
rect -3400 -12680 -1180 -12520
rect -1120 -12680 -1100 -12520
rect -3400 -12700 -1100 -12680
rect 400 -12520 1400 -12500
rect 400 -12680 420 -12520
rect 480 -12680 1400 -12520
rect 400 -12700 1400 -12680
rect -3400 -13120 -1300 -13100
rect -3400 -13280 -1380 -13120
rect -1320 -13280 -1300 -13120
rect -3400 -13300 -1300 -13280
rect 200 -13120 1400 -13100
rect 200 -13280 220 -13120
rect 280 -13280 1400 -13120
rect 200 -13300 1400 -13280
rect -3400 -13720 -1500 -13700
rect -3400 -13880 -1580 -13720
rect -1520 -13880 -1500 -13720
rect -3400 -13900 -1500 -13880
rect 0 -13720 1400 -13700
rect 0 -13880 20 -13720
rect 80 -13880 1400 -13720
rect 0 -13900 1400 -13880
rect -3400 -14320 -1700 -14300
rect -3400 -14480 -1780 -14320
rect -1720 -14480 -1700 -14320
rect -3400 -14500 -1700 -14480
rect -200 -14320 1400 -14300
rect -200 -14480 -180 -14320
rect -120 -14480 1400 -14320
rect -200 -14500 1400 -14480
rect 3600 -14800 3800 -8000
rect -3400 -14920 1400 -14900
rect -3400 -15080 -1980 -14920
rect -1920 -15080 1400 -14920
rect -3400 -15100 1400 -15080
rect 3000 -15000 3800 -14800
rect -3400 -15520 1400 -15500
rect -3400 -15680 -2180 -15520
rect -2120 -15680 1400 -15520
rect -3400 -15700 1400 -15680
rect -3400 -16120 1400 -16100
rect -3400 -16280 -2380 -16120
rect -2320 -16280 1400 -16120
rect -3400 -16300 1400 -16280
rect -3400 -17000 1200 -16600
rect -3400 -17320 1400 -17300
rect -3400 -17480 -2380 -17320
rect -2320 -17480 1400 -17320
rect -3400 -17500 1400 -17480
rect -3400 -17920 1400 -17900
rect -3400 -18080 -2180 -17920
rect -2120 -18080 1400 -17920
rect -3400 -18100 1400 -18080
rect -1220 -18500 -1100 -18480
rect -3400 -18520 1400 -18500
rect -3400 -18680 -1980 -18520
rect -1920 -18680 1400 -18520
rect -3400 -18700 1400 -18680
rect 3000 -18600 3200 -15000
rect 3600 -18600 3800 -15000
rect 3000 -18800 3800 -18600
rect -3400 -19120 1400 -19100
rect -3400 -19280 -1780 -19120
rect -1720 -19280 1400 -19120
rect -3400 -19300 1400 -19280
rect -3400 -19720 -1500 -19700
rect -3400 -19880 -1580 -19720
rect -1520 -19880 -1500 -19720
rect -3400 -19900 -1500 -19880
rect 0 -19720 1400 -19700
rect 0 -19880 20 -19720
rect 80 -19880 1400 -19720
rect 0 -19900 1400 -19880
rect -3400 -20320 -1300 -20300
rect -3400 -20480 -1380 -20320
rect -1320 -20480 -1300 -20320
rect -3400 -20500 -1300 -20480
rect 200 -20320 1400 -20300
rect 200 -20480 220 -20320
rect 280 -20480 1400 -20320
rect 200 -20500 1400 -20480
rect -3400 -20920 -1100 -20900
rect -3400 -21080 -1180 -20920
rect -1120 -21080 -1100 -20920
rect -3400 -21100 -1100 -21080
rect 400 -20920 1400 -20900
rect 400 -21080 420 -20920
rect 480 -21080 1400 -20920
rect 400 -21100 1400 -21080
rect -3400 -21520 -900 -21500
rect -3400 -21680 -980 -21520
rect -920 -21680 -900 -21520
rect -3400 -21700 -900 -21680
rect 600 -21520 1400 -21500
rect 600 -21680 620 -21520
rect 680 -21680 1400 -21520
rect 600 -21700 1400 -21680
rect -6494 -22390 -6268 -21804
rect -4744 -22390 -4548 -21804
rect -6494 -22586 -4548 -22390
use AND  x1
timestamp 1769198914
transform 1 0 900 0 1 -1500
box 100 -6089 3189 900
use AND  x2
timestamp 1769198914
transform 1 0 900 0 -1 -10500
box 100 -6089 3189 900
use AND  x3
timestamp 1769198914
transform 1 0 900 0 1 -12300
box 100 -6089 3189 900
use AND  x4
timestamp 1769198914
transform 1 0 900 0 -1 -21300
box 100 -6089 3189 900
use LOGIC_INV  x9
timestamp 1769198914
transform 1 0 -2000 0 1 9200
box -400 -9700 8600 -5400
<< labels >>
flabel metal1 1000 -17000 1200 -16800 0 FreeSans 256 0 0 0 VSS
port 18 nsew
flabel metal1 1000 -800 1200 -600 0 FreeSans 256 0 0 0 VDD
port 17 nsew
flabel metal1 3800 -3400 4000 -3200 0 FreeSans 256 0 0 0 LOGICOUT_0_2
port 16 nsew
flabel metal1 3800 -14200 4000 -14000 0 FreeSans 256 0 0 0 LOGICOUT_0_6
port 14 nsew
flabel metal1 3800 -19600 4000 -19400 0 FreeSans 256 0 0 0 LOGICOUT_0_8
port 13 nsew
flabel metal1 -2700 2600 -2500 2800 0 FreeSans 256 0 0 0 LOGICIN_0_2
port 12 nsew
flabel metal1 -2900 1200 -2700 1400 0 FreeSans 256 0 0 0 LOGICIN_0_4
port 11 nsew
flabel metal1 -3200 1000 -3000 1200 0 FreeSans 256 0 0 0 LOGICIN_0_6
port 10 nsew
flabel metal1 -3500 800 -3300 1000 0 FreeSans 256 0 0 0 LOGICIN_0_8
port 8 nsew
flabel metal1 -3800 600 -3600 800 0 FreeSans 256 0 0 0 LOGICIN_1_0
port 7 nsew
flabel metal1 -3600 300 -3400 500 0 FreeSans 256 0 0 0 LOGICIN_1_2
port 6 nsew
flabel metal1 -3300 100 -3100 300 0 FreeSans 256 0 0 0 LOGICIN_1_4
port 5 nsew
flabel metal1 -3000 -100 -2800 100 0 FreeSans 256 0 0 0 LOGICIN_1_6
port 4 nsew
flabel metal1 4000 -8800 4200 -8600 0 FreeSans 256 0 0 0 LOGICOUT_0_4
port 15 nsew
rlabel metal1 6710 -6926 7574 -6274 1 VSS
port 18 n
<< end >>
